magic
tech sky130A
magscale 1 2
timestamp 1757877451
<< locali >>
rect 73 1401 1125 1407
rect 73 1367 79 1401
rect 1119 1367 1125 1401
rect 73 1291 1125 1367
rect 73 -1240 1125 -1164
rect 73 -1274 79 -1240
rect 1119 -1274 1125 -1240
rect 73 -1280 1125 -1274
<< viali >>
rect 79 1367 1119 1401
rect 79 -1274 1119 -1240
<< metal1 >>
rect 37 1401 1161 1407
rect 37 1367 79 1401
rect 1119 1367 1161 1401
rect 37 1361 1161 1367
rect 133 1142 179 1361
rect 133 1127 181 1142
rect 133 1121 236 1127
rect 133 1096 178 1121
rect 172 1069 178 1096
rect 230 1069 236 1121
rect 172 1063 236 1069
rect 488 1121 552 1127
rect 488 1069 494 1121
rect 546 1069 552 1121
rect 488 1063 552 1069
rect 804 1121 868 1127
rect 804 1069 810 1121
rect 862 1069 868 1121
rect 804 1063 868 1069
rect 330 415 394 421
rect 330 363 336 415
rect 388 363 394 415
rect 330 357 394 363
rect 646 415 710 421
rect 646 363 652 415
rect 704 363 710 415
rect 646 357 710 363
rect 962 415 1026 421
rect 962 363 968 415
rect 1020 388 1026 415
rect 1020 363 1065 388
rect 962 357 1065 363
rect 1017 342 1065 357
rect 260 78 306 301
rect 418 78 464 301
rect 576 78 622 301
rect 734 78 780 307
rect 892 78 938 301
rect 260 32 938 78
rect 260 -192 306 32
rect 418 -192 464 32
rect 576 -192 622 32
rect 734 -186 780 32
rect 892 -186 938 32
rect 1019 -224 1065 342
rect 1017 -239 1065 -224
rect 330 -245 394 -239
rect 330 -297 336 -245
rect 388 -297 394 -245
rect 330 -303 394 -297
rect 646 -245 710 -239
rect 646 -297 652 -245
rect 704 -297 710 -245
rect 646 -303 710 -297
rect 962 -245 1065 -239
rect 962 -297 968 -245
rect 1020 -270 1065 -245
rect 1020 -297 1026 -270
rect 962 -303 1026 -297
rect 172 -951 236 -945
rect 172 -978 178 -951
rect 133 -1003 178 -978
rect 230 -1003 236 -951
rect 133 -1009 236 -1003
rect 488 -951 552 -945
rect 488 -1003 494 -951
rect 546 -1003 552 -951
rect 488 -1009 552 -1003
rect 804 -951 868 -945
rect 804 -1003 810 -951
rect 862 -1003 868 -951
rect 804 -1009 868 -1003
rect 133 -1024 181 -1009
rect 133 -1234 179 -1024
rect 37 -1240 1161 -1234
rect 37 -1274 79 -1240
rect 1119 -1274 1161 -1240
rect 37 -1280 1161 -1274
<< via1 >>
rect 178 1069 230 1121
rect 494 1069 546 1121
rect 810 1069 862 1121
rect 336 363 388 415
rect 652 363 704 415
rect 968 363 1020 415
rect 336 -297 388 -245
rect 652 -297 704 -245
rect 968 -297 1020 -245
rect 178 -1003 230 -951
rect 494 -1003 546 -951
rect 810 -1003 862 -951
<< metal2 >>
rect 172 1121 236 1127
rect 172 1069 178 1121
rect 230 1118 236 1121
rect 488 1121 552 1127
rect 488 1118 494 1121
rect 230 1072 494 1118
rect 230 1069 236 1072
rect 172 1063 236 1069
rect 488 1069 494 1072
rect 546 1118 552 1121
rect 804 1121 868 1127
rect 804 1118 810 1121
rect 546 1072 810 1118
rect 546 1069 552 1072
rect 488 1063 552 1069
rect 804 1069 810 1072
rect 862 1069 868 1121
rect 804 1063 868 1069
rect 330 415 394 421
rect 330 363 336 415
rect 388 412 394 415
rect 646 415 710 421
rect 646 412 652 415
rect 388 366 652 412
rect 388 363 394 366
rect 330 357 394 363
rect 646 363 652 366
rect 704 412 710 415
rect 962 415 1026 421
rect 962 412 968 415
rect 704 366 968 412
rect 704 363 710 366
rect 646 357 710 363
rect 962 363 968 366
rect 1020 363 1026 415
rect 962 357 1026 363
rect 330 -245 394 -239
rect 330 -297 336 -245
rect 388 -248 394 -245
rect 646 -245 710 -239
rect 646 -248 652 -245
rect 388 -294 652 -248
rect 388 -297 394 -294
rect 330 -303 394 -297
rect 646 -297 652 -294
rect 704 -248 710 -245
rect 962 -245 1026 -239
rect 962 -248 968 -245
rect 704 -294 968 -248
rect 704 -297 710 -294
rect 646 -303 710 -297
rect 962 -297 968 -294
rect 1020 -297 1026 -245
rect 962 -303 1026 -297
rect 172 -951 236 -945
rect 172 -1003 178 -951
rect 230 -954 236 -951
rect 488 -951 552 -945
rect 488 -954 494 -951
rect 230 -1000 494 -954
rect 230 -1003 236 -1000
rect 172 -1009 236 -1003
rect 488 -1003 494 -1000
rect 546 -954 552 -951
rect 804 -951 868 -945
rect 804 -954 810 -951
rect 546 -1000 810 -954
rect 546 -1003 552 -1000
rect 488 -1009 552 -1003
rect 804 -1003 810 -1000
rect 862 -1003 868 -951
rect 804 -1009 868 -1003
use sky130_fd_pr__nfet_01v8_TEWFY7  sky130_fd_pr__nfet_01v8_TEWFY7_0
timestamp 1757858607
transform 1 0 599 0 1 -624
box -562 -610 562 610
use sky130_fd_pr__pfet_01v8_X45PJH  sky130_fd_pr__pfet_01v8_X45PJH_0
timestamp 1757858607
transform 1 0 599 0 1 742
box -562 -619 562 619
<< end >>
