** sch_path: /foss/designs/mixedsignal/xschem/4-to-1_analog_MUX.sch
.subckt 4-to-1_analog_MUX S1 S2 VDD GND I1 I2 OUT I3 I4
*.PININFO I1:I I2:I I3:I I4:I OUT:O S1:I S2:I VDD:I GND:I
x1 S1 S1bar GND VDD Inverter
x2 S2 S2bar GND VDD Inverter
XM9 net1 S2 OUT VDD sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=1
XM1 I1 S1 net1 VDD sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=1
XM2 I3 S1bar net1 VDD sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=1
XM5 I2 S1 net2 VDD sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=1
XM7 I4 S1bar net2 VDD sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=1
XM11 net2 S2bar OUT VDD sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=1
XM3 I1 S1bar net1 GND sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM4 I3 S1 net1 GND sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM10 net1 S2bar OUT GND sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM6 I2 S1bar net2 GND sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM8 I4 S1 net2 GND sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM12 net2 S2 OUT GND sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
.ends

* expanding   symbol:  Inverter.sym # of pins=4
** sym_path: /foss/designs/mixedsignal/xschem/Inverter.sym
** sch_path: /foss/designs/mixedsignal/xschem/Inverter.sch
.subckt Inverter Vin Vout GND VDD
*.PININFO Vout:O Vin:I VDD:I GND:I
XM1 Vout Vin VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=1
XM2 Vout Vin GND GND sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
.ends

.end
