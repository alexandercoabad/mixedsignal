magic
tech sky130A
magscale 1 2
timestamp 1757874219
<< nwell >>
rect -712 -863 1656 -225
rect -712 -3153 1656 -2515
<< locali >>
rect -34 -185 1570 -179
rect -34 -219 -28 -185
rect 1564 -219 1570 -185
rect -34 -295 1570 -219
rect -84 -1626 1620 -1550
rect -84 -1660 -78 -1626
rect 1614 -1660 1620 -1626
rect -84 -1718 1620 -1660
rect -84 -1752 -78 -1718
rect 1614 -1752 1620 -1718
rect -84 -1828 1620 -1752
rect -34 -3159 1570 -3083
rect -34 -3193 -28 -3159
rect 1564 -3193 1570 -3159
rect -34 -3199 1570 -3193
<< viali >>
rect -28 -219 1564 -185
rect -78 -1660 1614 -1626
rect -78 -1752 1614 -1718
rect -28 -3193 1564 -3159
<< metal1 >>
rect -152 -176 -88 -170
rect -152 -179 -146 -176
rect -712 -225 -146 -179
rect -152 -228 -146 -225
rect -94 -179 -88 -176
rect -94 -185 1656 -179
rect -94 -219 -28 -185
rect 1564 -219 1656 -185
rect -94 -225 1656 -219
rect -94 -228 -88 -225
rect -152 -234 -88 -228
rect 657 -574 721 -568
rect 657 -598 663 -574
rect -24 -644 74 -598
rect 278 -626 663 -598
rect 715 -626 721 -574
rect 1249 -574 1313 -568
rect 1249 -598 1255 -574
rect 278 -632 721 -626
rect 278 -644 666 -632
rect 870 -644 968 -598
rect -448 -682 -384 -676
rect -448 -734 -442 -682
rect -390 -734 -384 -682
rect -448 -740 -384 -734
rect -439 -1178 -393 -740
rect -271 -1124 -207 -1118
rect -271 -1176 -265 -1124
rect -213 -1176 -207 -1124
rect -271 -1182 -207 -1176
rect -24 -1210 22 -644
rect 144 -682 208 -676
rect 144 -685 150 -682
rect 130 -731 150 -685
rect 144 -734 150 -731
rect 202 -685 208 -682
rect 202 -734 263 -685
rect 144 -740 263 -734
rect 97 -860 161 -854
rect 97 -912 103 -860
rect 155 -912 161 -860
rect 97 -918 161 -912
rect 106 -1118 152 -918
rect 217 -945 263 -740
rect 208 -951 272 -945
rect 208 -1003 214 -951
rect 266 -1003 272 -951
rect 208 -1009 272 -1003
rect 97 -1124 161 -1118
rect 97 -1132 103 -1124
rect 80 -1176 103 -1132
rect 155 -1132 161 -1124
rect 155 -1176 272 -1132
rect 80 -1178 272 -1176
rect 97 -1182 161 -1178
rect 330 -1210 376 -644
rect 568 -1210 614 -644
rect 681 -731 814 -685
rect 681 -854 727 -731
rect 672 -860 736 -854
rect 672 -912 678 -860
rect 730 -912 736 -860
rect 672 -918 736 -912
rect 783 -951 847 -945
rect 783 -1003 789 -951
rect 841 -1003 847 -951
rect 783 -1009 847 -1003
rect 792 -1178 838 -1009
rect 922 -1210 968 -644
rect -24 -1256 24 -1210
rect 328 -1222 616 -1210
rect 328 -1228 671 -1222
rect 328 -1256 613 -1228
rect 607 -1280 613 -1256
rect 665 -1280 671 -1228
rect 920 -1256 968 -1210
rect 1160 -626 1255 -598
rect 1307 -626 1313 -574
rect 1551 -595 1615 -589
rect 1551 -598 1557 -595
rect 1160 -632 1313 -626
rect 1160 -644 1258 -632
rect 1462 -644 1557 -598
rect 1160 -1210 1206 -644
rect 1551 -647 1557 -644
rect 1609 -647 1615 -595
rect 1551 -653 1615 -647
rect 1392 -682 1456 -676
rect 1392 -685 1398 -682
rect 1314 -731 1398 -685
rect 1392 -734 1398 -731
rect 1450 -734 1456 -682
rect 1392 -740 1456 -734
rect 1551 -1207 1615 -1201
rect 1551 -1210 1557 -1207
rect 1160 -1222 1208 -1210
rect 1160 -1228 1263 -1222
rect 1160 -1256 1205 -1228
rect 607 -1286 671 -1280
rect 1199 -1280 1205 -1256
rect 1257 -1280 1263 -1228
rect 1512 -1256 1557 -1210
rect 1551 -1259 1557 -1256
rect 1609 -1259 1615 -1207
rect 1551 -1265 1615 -1259
rect 1199 -1286 1263 -1280
rect 144 -1439 208 -1433
rect 144 -1491 150 -1439
rect 202 -1491 208 -1439
rect 144 -1497 208 -1491
rect 736 -1439 800 -1433
rect 736 -1491 742 -1439
rect 794 -1491 800 -1439
rect 736 -1497 800 -1491
rect 1264 -1444 1328 -1438
rect 1264 -1496 1270 -1444
rect 1322 -1496 1328 -1444
rect 1264 -1502 1328 -1496
rect -712 -1626 1656 -1620
rect -712 -1660 -78 -1626
rect 1614 -1660 1656 -1626
rect -712 -1718 1656 -1660
rect -712 -1752 -78 -1718
rect 1614 -1752 1656 -1718
rect -712 -1758 1656 -1752
rect 144 -1887 208 -1881
rect 144 -1939 150 -1887
rect 202 -1939 208 -1887
rect 144 -1945 208 -1939
rect 736 -1887 800 -1881
rect 736 -1939 742 -1887
rect 794 -1939 800 -1887
rect 736 -1945 800 -1939
rect 1392 -1883 1456 -1877
rect 1392 -1935 1398 -1883
rect 1450 -1935 1456 -1883
rect 1392 -1941 1456 -1935
rect 607 -2098 671 -2092
rect 607 -2122 613 -2098
rect -24 -2168 24 -2122
rect 328 -2150 613 -2122
rect 665 -2150 671 -2098
rect 1199 -2098 1263 -2092
rect 1199 -2122 1205 -2098
rect 328 -2156 671 -2150
rect 328 -2168 616 -2156
rect 920 -2168 968 -2122
rect -448 -2243 -384 -2237
rect -448 -2295 -442 -2243
rect -390 -2295 -384 -2243
rect -448 -2301 -384 -2295
rect -271 -2598 -207 -2592
rect -271 -2650 -265 -2598
rect -213 -2650 -207 -2598
rect -271 -2656 -207 -2650
rect -24 -2734 22 -2168
rect 106 -2460 152 -2200
rect 208 -2375 272 -2369
rect 208 -2427 214 -2375
rect 266 -2427 272 -2375
rect 208 -2433 272 -2427
rect 97 -2466 161 -2460
rect 97 -2518 103 -2466
rect 155 -2518 161 -2466
rect 97 -2524 161 -2518
rect 217 -2647 263 -2433
rect 130 -2693 263 -2647
rect 330 -2734 376 -2168
rect 568 -2734 614 -2168
rect 792 -2369 838 -2200
rect 783 -2375 847 -2369
rect 783 -2427 789 -2375
rect 841 -2427 847 -2375
rect 783 -2433 847 -2427
rect 672 -2466 736 -2460
rect 672 -2518 678 -2466
rect 730 -2518 736 -2466
rect 672 -2524 736 -2518
rect 681 -2647 727 -2524
rect 681 -2693 814 -2647
rect 922 -2734 968 -2168
rect -24 -2780 74 -2734
rect 278 -2746 666 -2734
rect 278 -2752 721 -2746
rect 278 -2780 663 -2752
rect 657 -2804 663 -2780
rect 715 -2804 721 -2752
rect 870 -2780 968 -2734
rect 1160 -2150 1205 -2122
rect 1257 -2150 1263 -2098
rect 1551 -2119 1615 -2113
rect 1551 -2122 1557 -2119
rect 1160 -2156 1263 -2150
rect 1160 -2168 1208 -2156
rect 1512 -2168 1557 -2122
rect 1160 -2734 1206 -2168
rect 1551 -2171 1557 -2168
rect 1609 -2171 1615 -2119
rect 1551 -2177 1615 -2171
rect 1264 -2644 1328 -2638
rect 1264 -2696 1270 -2644
rect 1322 -2647 1328 -2644
rect 1322 -2693 1406 -2647
rect 1322 -2696 1328 -2693
rect 1264 -2702 1328 -2696
rect 1551 -2731 1615 -2725
rect 1551 -2734 1557 -2731
rect 1160 -2746 1258 -2734
rect 1160 -2752 1313 -2746
rect 1160 -2780 1255 -2752
rect 657 -2810 721 -2804
rect 1249 -2804 1255 -2780
rect 1307 -2804 1313 -2752
rect 1462 -2780 1557 -2734
rect 1551 -2783 1557 -2780
rect 1609 -2783 1615 -2731
rect 1551 -2789 1615 -2783
rect 1249 -2810 1313 -2804
rect -152 -3150 -88 -3144
rect -152 -3202 -146 -3150
rect -94 -3153 -88 -3150
rect -94 -3159 1656 -3153
rect -94 -3193 -28 -3159
rect 1564 -3193 1656 -3159
rect -94 -3199 1656 -3193
rect -94 -3202 -88 -3199
rect -152 -3208 -88 -3202
<< via1 >>
rect -146 -228 -94 -176
rect 663 -626 715 -574
rect -442 -734 -390 -682
rect -265 -1176 -213 -1124
rect 150 -734 202 -682
rect 103 -912 155 -860
rect 214 -1003 266 -951
rect 103 -1176 155 -1124
rect 678 -912 730 -860
rect 789 -1003 841 -951
rect 613 -1280 665 -1228
rect 1255 -626 1307 -574
rect 1557 -647 1609 -595
rect 1398 -734 1450 -682
rect 1205 -1280 1257 -1228
rect 1557 -1259 1609 -1207
rect 150 -1491 202 -1439
rect 742 -1491 794 -1439
rect 1270 -1496 1322 -1444
rect 150 -1939 202 -1887
rect 742 -1939 794 -1887
rect 1398 -1935 1450 -1883
rect 613 -2150 665 -2098
rect -442 -2295 -390 -2243
rect -265 -2650 -213 -2598
rect 214 -2427 266 -2375
rect 103 -2518 155 -2466
rect 789 -2427 841 -2375
rect 678 -2518 730 -2466
rect 663 -2804 715 -2752
rect 1205 -2150 1257 -2098
rect 1557 -2171 1609 -2119
rect 1270 -2696 1322 -2644
rect 1255 -2804 1307 -2752
rect 1557 -2783 1609 -2731
rect -146 -3202 -94 -3150
<< metal2 >>
rect -157 -174 -83 -165
rect -157 -230 -148 -174
rect -92 -230 -83 -174
rect -157 -239 -83 -230
rect 657 -574 721 -568
rect 657 -626 663 -574
rect 715 -577 721 -574
rect 1249 -574 1313 -568
rect 1249 -577 1255 -574
rect 715 -623 1255 -577
rect 715 -626 721 -623
rect 657 -632 721 -626
rect 1249 -626 1255 -623
rect 1307 -626 1313 -574
rect 1249 -632 1313 -626
rect 1546 -593 1620 -584
rect 1546 -649 1555 -593
rect 1611 -649 1620 -593
rect 1546 -658 1620 -649
rect -448 -682 -384 -676
rect -448 -685 -442 -682
rect -462 -731 -442 -685
rect -448 -734 -442 -731
rect -390 -685 -384 -682
rect 144 -682 208 -676
rect 144 -685 150 -682
rect -390 -731 150 -685
rect -390 -734 -384 -731
rect -448 -740 -384 -734
rect 144 -734 150 -731
rect 202 -685 208 -682
rect 1387 -680 1461 -671
rect 202 -731 222 -685
rect 202 -734 208 -731
rect 144 -740 208 -734
rect 1387 -736 1396 -680
rect 1452 -736 1461 -680
rect 1387 -745 1461 -736
rect 97 -860 161 -854
rect 97 -912 103 -860
rect 155 -863 161 -860
rect 672 -860 736 -854
rect 672 -863 678 -860
rect 155 -909 678 -863
rect 155 -912 161 -909
rect 97 -918 161 -912
rect 672 -912 678 -909
rect 730 -912 736 -860
rect 672 -918 736 -912
rect 208 -951 272 -945
rect 208 -1003 214 -951
rect 266 -954 272 -951
rect 783 -951 847 -945
rect 783 -954 789 -951
rect 266 -1000 789 -954
rect 266 -1003 272 -1000
rect 208 -1009 272 -1003
rect 783 -1003 789 -1000
rect 841 -1003 847 -951
rect 783 -1009 847 -1003
rect -271 -1124 -207 -1118
rect -271 -1176 -265 -1124
rect -213 -1127 -207 -1124
rect 97 -1124 161 -1118
rect 97 -1127 103 -1124
rect -213 -1173 103 -1127
rect -213 -1176 -207 -1173
rect -271 -1182 -207 -1176
rect 97 -1176 103 -1173
rect 155 -1176 161 -1124
rect 97 -1182 161 -1176
rect 1546 -1205 1620 -1196
rect 607 -1228 671 -1222
rect 607 -1280 613 -1228
rect 665 -1231 671 -1228
rect 1199 -1228 1263 -1222
rect 1199 -1231 1205 -1228
rect 665 -1277 1205 -1231
rect 665 -1280 671 -1277
rect 607 -1286 671 -1280
rect 1199 -1280 1205 -1277
rect 1257 -1280 1263 -1228
rect 1546 -1261 1555 -1205
rect 1611 -1261 1620 -1205
rect 1546 -1270 1620 -1261
rect 1199 -1286 1263 -1280
rect 144 -1439 208 -1433
rect 144 -1491 150 -1439
rect 202 -1491 208 -1439
rect 144 -1497 208 -1491
rect 736 -1439 800 -1433
rect 736 -1491 742 -1439
rect 794 -1491 800 -1439
rect 736 -1497 800 -1491
rect 1259 -1442 1333 -1433
rect 153 -1881 199 -1497
rect 745 -1881 791 -1497
rect 1259 -1498 1268 -1442
rect 1324 -1498 1333 -1442
rect 1259 -1507 1333 -1498
rect 1387 -1881 1461 -1872
rect 144 -1887 208 -1881
rect 144 -1939 150 -1887
rect 202 -1939 208 -1887
rect 144 -1945 208 -1939
rect 736 -1887 800 -1881
rect 736 -1939 742 -1887
rect 794 -1939 800 -1887
rect 736 -1945 800 -1939
rect 1387 -1937 1396 -1881
rect 1452 -1937 1461 -1881
rect 1387 -1946 1461 -1937
rect 607 -2098 671 -2092
rect 607 -2150 613 -2098
rect 665 -2101 671 -2098
rect 1199 -2098 1263 -2092
rect 1199 -2101 1205 -2098
rect 665 -2147 1205 -2101
rect 665 -2150 671 -2147
rect 607 -2156 671 -2150
rect 1199 -2150 1205 -2147
rect 1257 -2150 1263 -2098
rect 1199 -2156 1263 -2150
rect 1546 -2117 1620 -2108
rect 1546 -2173 1555 -2117
rect 1611 -2173 1620 -2117
rect 1546 -2182 1620 -2173
rect -448 -2243 -384 -2237
rect -448 -2295 -442 -2243
rect -390 -2246 -384 -2243
rect 1387 -2241 1461 -2232
rect 1387 -2246 1396 -2241
rect -390 -2292 1396 -2246
rect -390 -2295 -384 -2292
rect -448 -2301 -384 -2295
rect 1387 -2297 1396 -2292
rect 1452 -2297 1461 -2241
rect 1387 -2306 1461 -2297
rect 208 -2375 272 -2369
rect 208 -2427 214 -2375
rect 266 -2378 272 -2375
rect 783 -2375 847 -2369
rect 783 -2378 789 -2375
rect 266 -2424 789 -2378
rect 266 -2427 272 -2424
rect 208 -2433 272 -2427
rect 783 -2427 789 -2424
rect 841 -2427 847 -2375
rect 783 -2433 847 -2427
rect 97 -2466 161 -2460
rect 97 -2518 103 -2466
rect 155 -2469 161 -2466
rect 672 -2466 736 -2460
rect 672 -2469 678 -2466
rect 155 -2515 678 -2469
rect 155 -2518 161 -2515
rect 97 -2524 161 -2518
rect 672 -2518 678 -2515
rect 730 -2518 736 -2466
rect 672 -2524 736 -2518
rect -271 -2598 -207 -2592
rect -271 -2650 -265 -2598
rect -213 -2601 -207 -2598
rect 1259 -2596 1333 -2587
rect 1259 -2601 1268 -2596
rect -213 -2647 1268 -2601
rect -213 -2650 -207 -2647
rect -271 -2656 -207 -2650
rect 1259 -2698 1268 -2647
rect 1324 -2698 1333 -2596
rect 1259 -2707 1333 -2698
rect 1546 -2729 1620 -2720
rect 657 -2752 721 -2746
rect 657 -2804 663 -2752
rect 715 -2755 721 -2752
rect 1249 -2752 1313 -2746
rect 1249 -2755 1255 -2752
rect 715 -2801 1255 -2755
rect 715 -2804 721 -2801
rect 657 -2810 721 -2804
rect 1249 -2804 1255 -2801
rect 1307 -2804 1313 -2752
rect 1546 -2785 1555 -2729
rect 1611 -2785 1620 -2729
rect 1546 -2794 1620 -2785
rect 1249 -2810 1313 -2804
rect -157 -3148 -83 -3139
rect -157 -3204 -148 -3148
rect -92 -3204 -83 -3148
rect -157 -3213 -83 -3204
<< via2 >>
rect -148 -176 -92 -174
rect -148 -228 -146 -176
rect -146 -228 -94 -176
rect -94 -228 -92 -176
rect -148 -230 -92 -228
rect 1555 -595 1611 -593
rect 1555 -647 1557 -595
rect 1557 -647 1609 -595
rect 1609 -647 1611 -595
rect 1555 -649 1611 -647
rect 1396 -682 1452 -680
rect 1396 -734 1398 -682
rect 1398 -734 1450 -682
rect 1450 -734 1452 -682
rect 1396 -736 1452 -734
rect 1555 -1207 1611 -1205
rect 1555 -1259 1557 -1207
rect 1557 -1259 1609 -1207
rect 1609 -1259 1611 -1207
rect 1555 -1261 1611 -1259
rect 1268 -1444 1324 -1442
rect 1268 -1496 1270 -1444
rect 1270 -1496 1322 -1444
rect 1322 -1496 1324 -1444
rect 1268 -1498 1324 -1496
rect 1396 -1883 1452 -1881
rect 1396 -1935 1398 -1883
rect 1398 -1935 1450 -1883
rect 1450 -1935 1452 -1883
rect 1396 -1937 1452 -1935
rect 1555 -2119 1611 -2117
rect 1555 -2171 1557 -2119
rect 1557 -2171 1609 -2119
rect 1609 -2171 1611 -2119
rect 1555 -2173 1611 -2171
rect 1396 -2297 1452 -2241
rect 1268 -2644 1324 -2596
rect 1268 -2696 1270 -2644
rect 1270 -2696 1322 -2644
rect 1322 -2696 1324 -2644
rect 1268 -2698 1324 -2696
rect 1555 -2731 1611 -2729
rect 1555 -2783 1557 -2731
rect 1557 -2783 1609 -2731
rect 1609 -2783 1611 -2731
rect 1555 -2785 1611 -2783
rect -148 -3150 -92 -3148
rect -148 -3202 -146 -3150
rect -146 -3202 -94 -3150
rect -94 -3202 -92 -3150
rect -148 -3204 -92 -3202
<< metal3 >>
rect -153 -174 -87 -169
rect -153 -230 -148 -174
rect -92 -230 -87 -174
rect -153 -235 -87 -230
rect -150 -3143 -90 -235
rect 1550 -593 1616 -588
rect 1550 -649 1555 -593
rect 1611 -649 1616 -593
rect 1550 -654 1616 -649
rect 1391 -680 1457 -675
rect 1391 -736 1396 -680
rect 1452 -736 1457 -680
rect 1391 -741 1457 -736
rect 1263 -1442 1329 -1437
rect 1263 -1498 1268 -1442
rect 1324 -1498 1329 -1442
rect 1263 -1503 1329 -1498
rect 1266 -2591 1326 -1503
rect 1394 -1876 1454 -741
rect 1553 -1200 1613 -654
rect 1550 -1205 1616 -1200
rect 1550 -1261 1555 -1205
rect 1611 -1261 1616 -1205
rect 1550 -1266 1616 -1261
rect 1391 -1881 1457 -1876
rect 1391 -1937 1396 -1881
rect 1452 -1937 1457 -1881
rect 1391 -1942 1457 -1937
rect 1394 -2236 1454 -1942
rect 1553 -2112 1613 -1266
rect 1550 -2117 1616 -2112
rect 1550 -2173 1555 -2117
rect 1611 -2173 1616 -2117
rect 1550 -2178 1616 -2173
rect 1391 -2241 1457 -2236
rect 1391 -2297 1396 -2241
rect 1452 -2297 1457 -2241
rect 1391 -2302 1457 -2297
rect 1263 -2596 1329 -2591
rect 1263 -2698 1268 -2596
rect 1324 -2698 1329 -2596
rect 1263 -2703 1329 -2698
rect 1553 -2724 1613 -2178
rect 1550 -2729 1616 -2724
rect 1550 -2785 1555 -2729
rect 1611 -2785 1616 -2729
rect 1550 -2790 1616 -2785
rect -153 -3148 -87 -3143
rect -153 -3204 -148 -3148
rect -92 -3204 -87 -3148
rect -153 -3209 -87 -3204
use Inverter  Inverter_0
timestamp 1757874219
transform 1 0 -2007 0 -1 -2731
box 1295 -1019 1887 468
use Inverter  Inverter_1
timestamp 1757874219
transform 1 0 -2007 0 1 -647
box 1295 -1019 1887 468
use sky130_fd_pr__nfet_01v8_JZTGL9  sky130_fd_pr__nfet_01v8_JZTGL9_0
timestamp 1757863532
transform 1 0 176 0 1 -1310
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_JZTGL9  sky130_fd_pr__nfet_01v8_JZTGL9_1
timestamp 1757863532
transform 1 0 768 0 -1 -2068
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_JZTGL9  sky130_fd_pr__nfet_01v8_JZTGL9_2
timestamp 1757863532
transform 1 0 176 0 -1 -2068
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_JZTGL9  sky130_fd_pr__nfet_01v8_JZTGL9_3
timestamp 1757863532
transform 1 0 1360 0 1 -1310
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_JZTGL9  sky130_fd_pr__nfet_01v8_JZTGL9_4
timestamp 1757863532
transform 1 0 768 0 1 -1310
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_JZTGL9  sky130_fd_pr__nfet_01v8_JZTGL9_5
timestamp 1757863532
transform 1 0 1360 0 -1 -2068
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_U6BDKB  sky130_fd_pr__pfet_01v8_U6BDKB_0
timestamp 1757863532
transform 1 0 1360 0 1 -544
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_U6BDKB  sky130_fd_pr__pfet_01v8_U6BDKB_1
timestamp 1757863532
transform 1 0 768 0 -1 -2834
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_U6BDKB  sky130_fd_pr__pfet_01v8_U6BDKB_2
timestamp 1757863532
transform 1 0 176 0 -1 -2834
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_U6BDKB  sky130_fd_pr__pfet_01v8_U6BDKB_3
timestamp 1757863532
transform 1 0 176 0 1 -544
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_U6BDKB  sky130_fd_pr__pfet_01v8_U6BDKB_4
timestamp 1757863532
transform 1 0 768 0 1 -544
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_U6BDKB  sky130_fd_pr__pfet_01v8_U6BDKB_5
timestamp 1757863532
transform 1 0 1360 0 -1 -2834
box -246 -319 246 319
<< labels >>
flabel metal1 922 -1256 968 -598 0 FreeSans 160 0 0 0 I3
port 3 nsew
flabel metal1 -24 -2780 22 -2122 0 FreeSans 160 0 0 0 I2
port 2 nsew
flabel metal1 922 -2780 968 -2122 0 FreeSans 160 0 0 0 I4
port 4 nsew
flabel metal3 1266 -2642 1326 -1498 0 FreeSans 160 90 0 0 S2bar
flabel metal1 -120 -1758 1656 -1620 0 FreeSans 320 0 0 0 GND
port 0 nsew
flabel metal1 -439 -1178 -393 -685 0 FreeSans 160 0 0 0 S1
port 5 nsew
flabel metal1 -439 -2301 -393 -2295 0 FreeSans 160 0 0 0 S2
port 6 nsew
flabel metal3 1394 -1881 1454 -736 0 FreeSans 160 90 0 0 S2
flabel metal1 -24 -1256 22 -598 0 FreeSans 160 0 0 0 I1
port 1 nsew
flabel metal1 -712 -225 1656 -179 0 FreeSans 160 0 0 0 VDD
port 7 nsew
flabel metal3 1553 -2783 1613 -595 0 FreeSans 160 90 0 0 OUT
port 9 nsew
<< end >>
