magic
tech sky130A
magscale 1 2
timestamp 1757870375
<< pwell >>
rect -739 -1442 739 1442
<< psubdiff >>
rect -703 1372 -607 1406
rect 607 1372 703 1406
rect -703 1310 -669 1372
rect 669 1310 703 1372
rect -703 -1372 -669 -1310
rect 669 -1372 703 -1310
rect -703 -1406 -607 -1372
rect 607 -1406 703 -1372
<< psubdiffcont >>
rect -607 1372 607 1406
rect -703 -1310 -669 1310
rect 669 -1310 703 1310
rect -607 -1406 607 -1372
<< xpolycontact >>
rect -573 844 573 1276
rect -573 -1276 573 -844
<< xpolyres >>
rect -573 -844 573 844
<< locali >>
rect -703 1372 -607 1406
rect 607 1372 703 1406
rect -703 1310 -669 1372
rect 669 1310 703 1372
rect -703 -1372 -669 -1310
rect 669 -1372 703 -1310
rect -703 -1406 -607 -1372
rect 607 -1406 703 -1372
<< viali >>
rect -557 861 557 1258
rect -557 -1258 557 -861
<< metal1 >>
rect -569 1258 569 1264
rect -569 861 -557 1258
rect 557 861 569 1258
rect -569 855 569 861
rect -569 -861 569 -855
rect -569 -1258 -557 -861
rect 557 -1258 569 -861
rect -569 -1264 569 -1258
<< properties >>
string FIXED_BBOX -686 -1389 686 1389
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 8.6 m 1 nx 1 wmin 5.730 lmin 0.50 class resistor rho 2000 val 3.067k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0 mult 1
<< end >>
