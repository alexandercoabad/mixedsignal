magic
tech sky130A
magscale 1 2
timestamp 1757870243
<< checkpaint >>
rect 6047 57453 10045 172159
rect 6047 17412 12895 57453
rect 4622 2202 12895 17412
rect 882 -266 12895 2202
rect -242 -3366 12895 -266
rect 3197 -3419 12895 -3366
rect 4622 -3472 12895 -3419
rect 6047 -3525 12895 -3472
rect 7472 -3578 12895 -3525
rect 8897 -3631 12895 -3578
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use 4-to-1_analog_MUX  x1
timestamp 1757868886
transform 1 0 2854 0 1 1107
box -712 -3213 1656 -165
use sky130_fd_pr__pfet_01v8_J9CDK9  XM3
timestamp 0
transform 1 0 509 0 1 -1754
box -562 -299 562 299
use sky130_fd_pr__nfet_01v8_TESQZT  XM4
timestamp 0
transform 1 0 1580 0 1 -1816
box -562 -290 562 290
use sky130_fd_pr__res_xhigh_po_5p73_PZF9TG  XR1
timestamp 0
transform 1 0 9471 0 1 -876
box -739 -1442 739 1442
use sky130_fd_pr__res_xhigh_po_5p73_UYUBYD  XR2
timestamp 0
transform 1 0 6621 0 1 6970
box -739 -9182 739 9182
use sky130_fd_pr__res_xhigh_po_5p73_PZF9TG  XR3
timestamp 0
transform 1 0 5196 0 1 -717
box -739 -1442 739 1442
use sky130_fd_pr__res_xhigh_po_5p73_86CYDR  XR4
timestamp 0
transform 1 0 8046 0 1 84317
box -739 -86582 739 86582
use sky130_fd_pr__res_xhigh_po_5p73_XKF2HR  XR5
timestamp 0
transform 1 0 10896 0 1 26911
box -739 -29282 739 29282
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 GND
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 S1
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 S2
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VIN
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VOUT
port 5 nsew
<< end >>
