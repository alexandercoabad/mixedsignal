magic
tech sky130A
magscale 1 2
timestamp 1757918270
<< locali >>
rect 15970 33511 30780 33545
rect 15970 30767 16106 33511
rect 15970 30627 30780 30767
rect 15970 27883 16106 30627
rect 15970 27743 30780 27883
rect 15970 24999 16106 27743
rect 15970 24859 30780 24999
rect 15970 22115 16106 24859
rect 15970 22082 30780 22115
rect 1262 22048 30780 22082
rect 15970 21975 30780 22048
rect 15970 20450 16106 21975
rect 1262 20310 16106 20450
rect 15970 19231 16106 20310
rect 15970 19091 30780 19231
rect 15970 18712 16106 19091
rect 1262 18572 16106 18712
rect 15970 16974 16106 18572
rect 1262 16834 16106 16974
rect 15970 16347 16106 16834
rect 15970 16207 30780 16347
rect 15970 15236 16106 16207
rect 1262 15096 16106 15236
rect 15970 13498 16106 15096
rect 1262 13463 16106 13498
rect 1262 13358 30780 13463
rect 15970 13323 30780 13358
rect 15970 11760 16106 13323
rect 1262 11620 16106 11760
rect 15970 10579 16106 11620
rect 15970 10439 30780 10579
rect 15970 10022 16106 10439
rect 1262 9882 16106 10022
rect 15970 8284 16106 9882
rect 1262 8144 16106 8284
rect 15970 7695 16106 8144
rect 15970 7555 30780 7695
rect 15970 6546 16106 7555
rect 1262 6406 16106 6546
rect 15970 4811 16106 6406
rect 15970 4808 30780 4811
rect 1262 4287 30780 4808
rect 1262 4098 20559 4287
rect 1262 4046 1744 4098
rect 1796 4046 20559 4098
rect 1262 3810 20559 4046
rect 1262 1054 2212 3810
rect 16862 3665 20559 3810
rect 16873 1054 18188 3665
rect 19539 2495 20559 3665
rect 22927 4264 30780 4287
rect 22927 3404 28884 4264
rect 22927 2495 25905 3404
rect 19529 2357 25905 2495
rect 1262 908 18188 1054
rect 19539 908 20559 2357
rect 1262 782 20559 908
rect 22927 782 25905 2357
rect 1262 771 25905 782
rect 27276 1530 28884 3404
rect 30008 1530 30780 4264
rect 1262 633 25899 771
rect 27276 633 30780 1530
rect 1262 405 30780 633
<< viali >>
rect 1744 4046 1796 4098
<< metal1 >>
rect 28971 4113 29035 4119
rect 1732 4098 1808 4110
rect 1732 4046 1744 4098
rect 1796 4046 1808 4098
rect 28971 4061 28977 4113
rect 29029 4061 29035 4113
rect 28971 4055 29035 4061
rect 1732 4034 1808 4046
rect 22184 3342 22248 3348
rect 22184 3290 22190 3342
rect 22242 3290 22248 3342
rect 22184 3284 22248 3290
rect 20823 3213 20887 3219
rect 20823 3161 20829 3213
rect 20881 3161 20887 3213
rect 20823 3155 20887 3161
rect 26556 3109 26620 3115
rect 26556 3057 26562 3109
rect 26614 3057 26620 3109
rect 26556 3051 26620 3057
rect 28629 3109 28693 3115
rect 28629 3057 28635 3109
rect 28687 3057 28693 3109
rect 28629 3051 28693 3057
rect 28638 2790 28684 3051
rect 28629 2784 28693 2790
rect 28629 2732 28635 2784
rect 28687 2732 28693 2784
rect 28629 2726 28693 2732
rect 29098 2784 29162 2790
rect 29098 2732 29104 2784
rect 29156 2732 29162 2784
rect 29098 2726 29162 2732
rect 29857 2784 29921 2790
rect 29857 2732 29863 2784
rect 29915 2732 29921 2784
rect 29857 2726 29921 2732
rect 20823 1716 20887 1722
rect 20823 1664 20829 1716
rect 20881 1664 20887 1716
rect 20823 1658 20887 1664
rect 21242 1717 21306 1723
rect 21242 1665 21248 1717
rect 21300 1665 21306 1717
rect 21242 1659 21306 1665
rect 22184 1708 22248 1714
rect 22184 1656 22190 1708
rect 22242 1656 22248 1708
rect 22184 1650 22248 1656
<< via1 >>
rect 1939 5110 1991 5162
rect 15241 5092 15293 5144
rect 17034 5109 17086 5161
rect 30426 5075 30478 5127
rect 1744 4046 1796 4098
rect 28977 4061 29029 4113
rect 19228 3290 19280 3342
rect 22190 3290 22242 3342
rect 20829 3161 20881 3213
rect 26562 3057 26614 3109
rect 28635 3057 28687 3109
rect 28635 2732 28687 2784
rect 29104 2732 29156 2784
rect 29863 2732 29915 2784
rect 20829 1664 20881 1716
rect 21248 1665 21300 1717
rect 22190 1656 22242 1708
rect 2865 1351 2917 1403
rect 16167 1350 16219 1402
rect 18834 1209 18886 1261
rect 26562 937 26614 989
<< metal2 >>
rect 20714 44218 20788 44227
rect 20714 44162 20723 44218
rect 20779 44213 20788 44218
rect 27103 44218 27177 44227
rect 27103 44213 27112 44218
rect 20779 44167 27112 44213
rect 20779 44162 20788 44167
rect 20714 44153 20788 44162
rect 27103 44162 27112 44167
rect 27168 44162 27177 44218
rect 27103 44153 27177 44162
rect 20909 43944 20983 43953
rect 20909 43888 20918 43944
rect 20974 43939 20983 43944
rect 27655 43944 27729 43953
rect 27655 43939 27664 43944
rect 20974 43893 27664 43939
rect 20974 43888 20983 43893
rect 20909 43879 20983 43888
rect 27655 43888 27664 43893
rect 27720 43888 27729 43944
rect 27655 43879 27729 43888
rect 1928 5164 2002 5173
rect 1928 5108 1937 5164
rect 1993 5108 2002 5164
rect 17023 5163 17097 5172
rect 1928 5099 2002 5108
rect 15230 5146 15304 5155
rect 15230 5090 15239 5146
rect 15295 5090 15304 5146
rect 17023 5107 17032 5163
rect 17088 5107 17097 5163
rect 17023 5098 17097 5107
rect 30415 5129 30489 5138
rect 15230 5081 15304 5090
rect 30415 5073 30424 5129
rect 30480 5073 30489 5129
rect 30415 5064 30489 5073
rect 1671 4512 1745 4521
rect 1671 4456 1680 4512
rect 1736 4507 1745 4512
rect 21114 4512 21188 4521
rect 21114 4507 21123 4512
rect 1736 4461 21123 4507
rect 1736 4456 1745 4461
rect 1671 4447 1745 4456
rect 21114 4456 21123 4461
rect 21179 4507 21188 4512
rect 28966 4512 29040 4521
rect 28966 4507 28975 4512
rect 21179 4461 28975 4507
rect 21179 4456 21188 4461
rect 21114 4447 21188 4456
rect 28966 4456 28975 4461
rect 29031 4456 29040 4512
rect 28966 4447 29040 4456
rect 15230 4231 15304 4240
rect 15230 4175 15239 4231
rect 15295 4226 15304 4231
rect 22179 4231 22253 4240
rect 22179 4226 22188 4231
rect 15295 4180 22188 4226
rect 15295 4175 15304 4180
rect 15230 4166 15304 4175
rect 22179 4175 22188 4180
rect 22244 4175 22253 4231
rect 22179 4166 22253 4175
rect 28966 4115 29040 4124
rect 1733 4100 1807 4109
rect 1733 4044 1742 4100
rect 1798 4044 1807 4100
rect 1733 4035 1807 4044
rect 17023 4078 17097 4087
rect 17023 4022 17032 4078
rect 17088 4073 17097 4078
rect 22817 4078 22891 4087
rect 22817 4073 22826 4078
rect 17088 4027 22826 4073
rect 17088 4022 17097 4027
rect 17023 4013 17097 4022
rect 22817 4022 22826 4027
rect 22882 4022 22891 4078
rect 28966 4059 28975 4115
rect 29031 4059 29040 4115
rect 28966 4050 29040 4059
rect 22817 4013 22891 4022
rect 19222 3342 19286 3348
rect 19222 3290 19228 3342
rect 19280 3339 19286 3342
rect 22184 3342 22248 3348
rect 22184 3339 22190 3342
rect 19280 3293 22190 3339
rect 19280 3290 19286 3293
rect 19222 3284 19286 3290
rect 22184 3290 22190 3293
rect 22242 3290 22248 3342
rect 22184 3284 22248 3290
rect 20714 3215 20788 3224
rect 20714 3159 20723 3215
rect 20779 3210 20788 3215
rect 20823 3213 20887 3219
rect 20823 3210 20829 3213
rect 20779 3164 20829 3210
rect 20779 3159 20788 3164
rect 20714 3150 20788 3159
rect 20823 3161 20829 3164
rect 20881 3161 20887 3213
rect 20823 3155 20887 3161
rect 22817 3111 22891 3120
rect 22817 3055 22826 3111
rect 22882 3106 22891 3111
rect 26556 3109 26620 3115
rect 26556 3106 26562 3109
rect 22882 3060 26562 3106
rect 22882 3055 22891 3060
rect 22817 3046 22891 3055
rect 26556 3057 26562 3060
rect 26614 3106 26620 3109
rect 28629 3109 28693 3115
rect 28629 3106 28635 3109
rect 26614 3060 28635 3106
rect 26614 3057 26620 3060
rect 26556 3051 26620 3057
rect 28629 3057 28635 3060
rect 28687 3057 28693 3109
rect 28629 3051 28693 3057
rect 28629 2784 28693 2790
rect 28629 2732 28635 2784
rect 28687 2781 28693 2784
rect 29098 2784 29162 2790
rect 29098 2781 29104 2784
rect 28687 2735 29104 2781
rect 28687 2732 28693 2735
rect 28629 2726 28693 2732
rect 29098 2732 29104 2735
rect 29156 2732 29162 2784
rect 29098 2726 29162 2732
rect 29857 2784 29921 2790
rect 29857 2732 29863 2784
rect 29915 2781 29921 2784
rect 30415 2786 30489 2795
rect 30415 2781 30424 2786
rect 29915 2735 30424 2781
rect 29915 2732 29921 2735
rect 29857 2726 29921 2732
rect 30415 2730 30424 2735
rect 30480 2730 30489 2786
rect 30415 2721 30489 2730
rect 20909 1722 20983 1727
rect 20823 1718 20983 1722
rect 20823 1716 20918 1718
rect 20823 1664 20829 1716
rect 20881 1664 20918 1716
rect 20823 1662 20918 1664
rect 20974 1662 20983 1718
rect 20823 1658 20983 1662
rect 20909 1653 20983 1658
rect 21237 1719 21311 1728
rect 21237 1663 21246 1719
rect 21302 1663 21311 1719
rect 21237 1654 21311 1663
rect 22179 1710 22253 1719
rect 22179 1654 22188 1710
rect 22244 1654 22253 1710
rect 22179 1645 22253 1654
rect 2854 1405 2928 1414
rect 2854 1349 2863 1405
rect 2919 1349 2928 1405
rect 2854 1340 2928 1349
rect 16156 1404 16230 1413
rect 16156 1348 16165 1404
rect 16221 1348 16230 1404
rect 16156 1339 16230 1348
rect 18823 1263 18897 1272
rect 18823 1207 18832 1263
rect 18888 1207 18897 1263
rect 18823 1198 18897 1207
rect 26551 991 26625 1000
rect 26551 935 26560 991
rect 26616 935 26625 991
rect 26551 926 26625 935
rect 16156 737 16230 746
rect 16156 681 16165 737
rect 16221 732 16230 737
rect 21237 737 21311 746
rect 21237 732 21246 737
rect 16221 686 21246 732
rect 16221 681 16230 686
rect 16156 672 16230 681
rect 21237 681 21246 686
rect 21302 681 21311 737
rect 21237 672 21311 681
rect 1928 391 2002 400
rect 1928 335 1937 391
rect 1993 386 2002 391
rect 2854 391 2928 400
rect 2854 386 2863 391
rect 1993 340 2863 386
rect 1993 335 2002 340
rect 1928 326 2002 335
rect 2854 335 2863 340
rect 2919 386 2928 391
rect 18823 391 18897 400
rect 18823 386 18832 391
rect 2919 340 18832 386
rect 2919 335 2928 340
rect 2854 326 2928 335
rect 18823 335 18832 340
rect 18888 386 18897 391
rect 30415 391 30489 400
rect 30415 386 30424 391
rect 18888 340 30424 386
rect 18888 335 18897 340
rect 18823 326 18897 335
rect 30415 335 30424 340
rect 30480 335 30489 391
rect 30415 326 30489 335
<< via2 >>
rect 20723 44162 20779 44218
rect 27112 44162 27168 44218
rect 20918 43888 20974 43944
rect 27664 43888 27720 43944
rect 1937 5162 1993 5164
rect 1937 5110 1939 5162
rect 1939 5110 1991 5162
rect 1991 5110 1993 5162
rect 1937 5108 1993 5110
rect 15239 5144 15295 5146
rect 15239 5092 15241 5144
rect 15241 5092 15293 5144
rect 15293 5092 15295 5144
rect 15239 5090 15295 5092
rect 17032 5161 17088 5163
rect 17032 5109 17034 5161
rect 17034 5109 17086 5161
rect 17086 5109 17088 5161
rect 17032 5107 17088 5109
rect 30424 5127 30480 5129
rect 30424 5075 30426 5127
rect 30426 5075 30478 5127
rect 30478 5075 30480 5127
rect 30424 5073 30480 5075
rect 1680 4456 1736 4512
rect 21123 4456 21179 4512
rect 28975 4456 29031 4512
rect 15239 4175 15295 4231
rect 22188 4175 22244 4231
rect 1742 4098 1798 4100
rect 1742 4046 1744 4098
rect 1744 4046 1796 4098
rect 1796 4046 1798 4098
rect 1742 4044 1798 4046
rect 17032 4022 17088 4078
rect 22826 4022 22882 4078
rect 28975 4113 29031 4115
rect 28975 4061 28977 4113
rect 28977 4061 29029 4113
rect 29029 4061 29031 4113
rect 28975 4059 29031 4061
rect 20723 3159 20779 3215
rect 22826 3055 22882 3111
rect 30424 2730 30480 2786
rect 20918 1662 20974 1718
rect 21246 1717 21302 1719
rect 21246 1665 21248 1717
rect 21248 1665 21300 1717
rect 21300 1665 21302 1717
rect 21246 1663 21302 1665
rect 22188 1708 22244 1710
rect 22188 1656 22190 1708
rect 22190 1656 22242 1708
rect 22242 1656 22244 1708
rect 22188 1654 22244 1656
rect 2863 1403 2919 1405
rect 2863 1351 2865 1403
rect 2865 1351 2917 1403
rect 2917 1351 2919 1403
rect 2863 1349 2919 1351
rect 16165 1402 16221 1404
rect 16165 1350 16167 1402
rect 16167 1350 16219 1402
rect 16219 1350 16221 1402
rect 16165 1348 16221 1350
rect 18832 1261 18888 1263
rect 18832 1209 18834 1261
rect 18834 1209 18886 1261
rect 18886 1209 18888 1261
rect 18832 1207 18888 1209
rect 26560 989 26616 991
rect 26560 937 26562 989
rect 26562 937 26614 989
rect 26614 937 26616 989
rect 26560 935 26616 937
rect 16165 681 16221 737
rect 21246 681 21302 737
rect 1937 335 1993 391
rect 2863 335 2919 391
rect 18832 335 18888 391
rect 30424 335 30480 391
<< metal3 >>
rect 27102 45005 27178 45011
rect 27102 44941 27108 45005
rect 27172 44941 27178 45005
rect 27102 44935 27178 44941
rect 27654 44997 27730 45003
rect 27110 44223 27170 44935
rect 27654 44933 27660 44997
rect 27724 44933 27730 44997
rect 27654 44927 27730 44933
rect 20718 44218 20784 44223
rect 20718 44162 20723 44218
rect 20779 44162 20784 44218
rect 20718 44157 20784 44162
rect 27107 44218 27173 44223
rect 27107 44162 27112 44218
rect 27168 44162 27173 44218
rect 27107 44157 27173 44162
rect 1932 5164 1998 5169
rect 1932 5108 1937 5164
rect 1993 5108 1998 5164
rect 17027 5163 17093 5168
rect 1932 5103 1998 5108
rect 15234 5146 15300 5151
rect 372 4534 484 4540
rect 372 4434 378 4534
rect 478 4514 484 4534
rect 1675 4514 1741 4517
rect 478 4512 1741 4514
rect 478 4456 1680 4512
rect 1736 4456 1741 4512
rect 478 4454 1741 4456
rect 478 4434 484 4454
rect 1675 4451 1741 4454
rect 372 4428 484 4434
rect 927 4122 1039 4128
rect 927 4022 933 4122
rect 1033 4102 1039 4122
rect 1737 4102 1803 4105
rect 1033 4100 1803 4102
rect 1033 4044 1742 4100
rect 1798 4044 1803 4100
rect 1033 4042 1803 4044
rect 1033 4022 1039 4042
rect 1737 4039 1803 4042
rect 927 4016 1039 4022
rect 1935 396 1995 5103
rect 15234 5090 15239 5146
rect 15295 5090 15300 5146
rect 17027 5107 17032 5163
rect 17088 5107 17093 5163
rect 17027 5102 17093 5107
rect 15234 5085 15300 5090
rect 15237 4236 15297 5085
rect 15234 4231 15300 4236
rect 15234 4175 15239 4231
rect 15295 4175 15300 4231
rect 15234 4170 15300 4175
rect 17030 4083 17090 5102
rect 17027 4078 17093 4083
rect 17027 4022 17032 4078
rect 17088 4022 17093 4078
rect 17027 4017 17093 4022
rect 20721 3220 20781 44157
rect 27662 43949 27722 44927
rect 20913 43944 20979 43949
rect 20913 43888 20918 43944
rect 20974 43888 20979 43944
rect 20913 43883 20979 43888
rect 27659 43944 27725 43949
rect 27659 43888 27664 43944
rect 27720 43888 27725 43944
rect 27659 43883 27725 43888
rect 20718 3215 20784 3220
rect 20718 3159 20723 3215
rect 20779 3159 20784 3215
rect 20718 3154 20784 3159
rect 20916 1723 20976 43883
rect 30419 5129 30485 5134
rect 30419 5073 30424 5129
rect 30480 5073 30485 5129
rect 30419 5068 30485 5073
rect 21118 4512 21184 4517
rect 21118 4456 21123 4512
rect 21179 4456 21184 4512
rect 21118 4451 21184 4456
rect 28970 4512 29036 4517
rect 28970 4456 28975 4512
rect 29031 4456 29036 4512
rect 28970 4451 29036 4456
rect 21121 3880 21181 4451
rect 22183 4231 22249 4236
rect 22183 4175 22188 4231
rect 22244 4175 22249 4231
rect 22183 4170 22249 4175
rect 20913 1718 20979 1723
rect 20913 1662 20918 1718
rect 20974 1662 20979 1718
rect 20913 1657 20979 1662
rect 21241 1719 21307 1724
rect 21241 1663 21246 1719
rect 21302 1663 21307 1719
rect 22186 1715 22246 4170
rect 28973 4120 29033 4451
rect 28970 4115 29036 4120
rect 22821 4078 22887 4083
rect 22821 4022 22826 4078
rect 22882 4022 22887 4078
rect 28970 4059 28975 4115
rect 29031 4059 29036 4115
rect 28970 4054 29036 4059
rect 22821 4017 22887 4022
rect 22824 3461 22884 4017
rect 22821 3111 22887 3116
rect 22821 3055 22826 3111
rect 22882 3055 22887 3111
rect 22821 3050 22887 3055
rect 30422 2791 30482 5068
rect 30419 2786 30485 2791
rect 30419 2730 30424 2786
rect 30480 2730 30485 2786
rect 30419 2725 30485 2730
rect 21241 1658 21307 1663
rect 22183 1710 22249 1715
rect 2858 1405 2924 1410
rect 2858 1349 2863 1405
rect 2919 1349 2924 1405
rect 2858 1344 2924 1349
rect 16160 1404 16226 1409
rect 16160 1348 16165 1404
rect 16221 1348 16226 1404
rect 2861 396 2921 1344
rect 16160 1343 16226 1348
rect 16163 742 16223 1343
rect 18827 1263 18893 1268
rect 18827 1207 18832 1263
rect 18888 1207 18893 1263
rect 18827 1202 18893 1207
rect 16160 737 16226 742
rect 16160 681 16165 737
rect 16221 681 16226 737
rect 16160 676 16226 681
rect 18830 396 18890 1202
rect 21244 742 21304 1658
rect 22183 1654 22188 1710
rect 22244 1654 22249 1710
rect 22183 1649 22249 1654
rect 26555 991 26621 996
rect 26555 935 26560 991
rect 26616 935 26621 991
rect 26555 930 26621 935
rect 21241 737 21307 742
rect 21241 681 21246 737
rect 21302 681 21307 737
rect 21241 676 21307 681
rect 1932 391 1998 396
rect 1932 335 1937 391
rect 1993 335 1998 391
rect 1932 330 1998 335
rect 2858 391 2924 396
rect 2858 335 2863 391
rect 2919 335 2924 391
rect 2858 330 2924 335
rect 18827 391 18893 396
rect 18827 335 18832 391
rect 18888 335 18893 391
rect 18827 330 18893 335
rect 26558 200 26618 930
rect 30422 396 30482 2725
rect 30419 391 30485 396
rect 30419 335 30424 391
rect 30480 335 30485 391
rect 30419 330 30485 335
rect 30422 200 30482 330
rect 26550 194 26626 200
rect 26550 130 26556 194
rect 26620 130 26626 194
rect 26550 124 26626 130
rect 30414 194 30490 200
rect 30414 130 30420 194
rect 30484 130 30490 194
rect 30414 124 30490 130
<< via3 >>
rect 27108 44941 27172 45005
rect 27660 44933 27724 44997
rect 378 4434 478 4534
rect 933 4022 1033 4122
rect 26556 130 26620 194
rect 30420 130 30484 194
<< metal4 >>
rect 27110 45006 27170 45152
rect 27107 45005 27173 45006
rect 27107 44941 27108 45005
rect 27172 44941 27173 45005
rect 27662 44998 27722 45152
rect 27107 44940 27173 44941
rect 27659 44997 27725 44998
rect 27659 44933 27660 44997
rect 27724 44933 27725 44997
rect 27659 44932 27725 44933
rect 200 4534 600 44152
rect 200 4434 378 4534
rect 478 4434 600 4534
rect 200 1000 600 4434
rect 800 4122 1200 44152
rect 800 4022 933 4122
rect 1033 4022 1200 4122
rect 800 1000 1200 4022
rect 26498 194 26678 200
rect 26498 130 26556 194
rect 26620 130 26678 194
rect 26498 0 26678 130
rect 30362 194 30542 200
rect 30362 130 30420 194
rect 30484 130 30542 194
rect 30362 0 30542 130
use 3k_res  3k_res_0
timestamp 1757918270
transform -1 0 27274 0 -1 3412
box -53 -53 1425 2831
use 3k_res  3k_res_1
timestamp 1757918270
transform 1 0 18174 0 1 904
box -53 -53 1425 2831
use 4-to-1_analog_MUX  4-to-1_analog_MUX_0
timestamp 1757918270
transform 1 0 21271 0 1 4115
box -712 -3213 1656 -165
use 30k_res  30k_res_0
timestamp 1757918270
transform -1 0 16847 0 1 1047
box -85 -51 14695 2833
use 100k_res  100k_res_1
timestamp 1757872436
transform -1 0 15919 0 1 4785
box -87 -47 14693 17333
use 300k_res  300k_res_1
timestamp 1757918270
transform -1 0 35651 0 1 -23932
box 4835 28673 19615 57513
use Inverter_base  Inverter_base_0
timestamp 1757877451
transform 1 0 28847 0 1 2703
box 37 -1280 1161 1407
<< labels >>
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal2 s 22882 3060 26562 3106 0 FreeSans 160 0 0 0 mux_in
<< properties >>
string (UNNAMED) gencell
string FIXED_BBOX 0 0 32200 45152
<< end >>
