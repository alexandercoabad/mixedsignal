magic
tech sky130A
magscale 1 2
timestamp 1740500291
<< nwell >>
rect 4762 8290 5464 12510
<< nmos >>
rect 5102 4050 5202 8050
<< pmos >>
rect 5102 8400 5202 12400
<< ndiff >>
rect 4882 8020 5102 8050
rect 4882 4080 4972 8020
rect 5012 4080 5102 8020
rect 4882 4050 5102 4080
rect 5202 8020 5422 8050
rect 5202 4080 5292 8020
rect 5332 4080 5422 8020
rect 5202 4050 5422 4080
<< pdiff >>
rect 4882 12370 5102 12400
rect 4882 8430 4972 12370
rect 5012 8430 5102 12370
rect 4882 8400 5102 8430
rect 5202 12370 5422 12400
rect 5202 8430 5292 12370
rect 5332 8430 5422 12370
rect 5202 8400 5422 8430
<< ndiffc >>
rect 4972 4080 5012 8020
rect 5292 4080 5332 8020
<< pdiffc >>
rect 4972 8430 5012 12370
rect 5292 8430 5332 12370
<< psubdiff >>
rect 4802 8020 4882 8050
rect 4802 4080 4822 8020
rect 4862 4080 4882 8020
rect 4802 4050 4882 4080
<< nsubdiff >>
rect 4802 12370 4882 12400
rect 4802 8430 4822 12370
rect 4862 8430 4882 12370
rect 4802 8400 4882 8430
<< psubdiffcont >>
rect 4822 4080 4862 8020
<< nsubdiffcont >>
rect 4822 8430 4862 12370
<< poly >>
rect 5102 12400 5202 12500
rect 5102 8290 5202 8400
rect 5022 8280 5202 8290
rect 5022 8240 5042 8280
rect 5082 8240 5202 8280
rect 5022 8230 5202 8240
rect 5102 8050 5202 8230
rect 5102 3950 5202 4050
<< polycont >>
rect 5042 8240 5082 8280
<< locali >>
rect 4802 12390 4842 12440
rect 4802 12370 5092 12390
rect 4802 8430 4822 12370
rect 4862 8430 4972 12370
rect 5012 8430 5092 12370
rect 4802 8410 5092 8430
rect 5212 12370 5422 12390
rect 5212 8430 5292 12370
rect 5332 8430 5422 12370
rect 5212 8290 5422 8430
rect 4742 8280 5102 8290
rect 4742 8240 4762 8280
rect 4802 8240 5042 8280
rect 5082 8240 5102 8280
rect 4742 8230 5102 8240
rect 5212 8280 5622 8290
rect 5212 8240 5562 8280
rect 5602 8240 5622 8280
rect 5212 8230 5622 8240
rect 4802 8020 5092 8040
rect 4802 4080 4822 8020
rect 4862 4080 4972 8020
rect 5012 4080 5092 8020
rect 4802 4060 5092 4080
rect 5212 8020 5422 8230
rect 5212 4080 5292 8020
rect 5332 4080 5422 8020
rect 5212 4060 5422 4080
rect 4802 4010 4842 4060
<< viali >>
rect 4800 12440 4842 12480
rect 4762 8240 4802 8280
rect 5562 8240 5602 8280
rect 4802 3970 4842 4010
<< metal1 >>
rect 4252 19130 5612 19200
rect 4500 12430 4520 12490
rect 4580 12480 5482 12490
rect 4580 12440 4800 12480
rect 4842 12440 5482 12480
rect 4580 12430 5482 12440
rect 3200 9870 3580 9940
rect 3200 8540 3350 9870
rect 3200 8430 3220 8540
rect 3330 8430 3350 8540
rect 3512 8290 3582 8890
rect 5542 8290 5612 19130
rect 5980 8290 6060 8300
rect 3512 8280 4822 8290
rect 3512 8240 4762 8280
rect 4802 8240 4822 8280
rect 3512 8230 4822 8240
rect 5540 8280 5990 8290
rect 5540 8240 5562 8280
rect 5602 8240 5990 8280
rect 5540 8230 5990 8240
rect 6050 8230 6060 8290
rect 5980 8220 6060 8230
rect 4430 4030 4530 4040
rect 4430 3950 4440 4030
rect 4520 4020 4530 4030
rect 4520 4010 5482 4020
rect 4520 3970 4802 4010
rect 4842 3970 5482 4010
rect 4520 3960 5482 3970
rect 4520 3950 4530 3960
rect 4430 3940 4530 3950
<< via1 >>
rect 4520 12430 4580 12490
rect 3220 8430 3330 8540
rect 5990 8230 6050 8290
rect 4440 3950 4520 4030
<< metal2 >>
rect 4310 12500 4410 12510
rect 4310 12420 4320 12500
rect 4400 12490 4410 12500
rect 4400 12430 4520 12490
rect 4580 12430 4590 12490
rect 4400 12420 4410 12430
rect 4310 12410 4410 12420
rect 3200 8540 3350 8550
rect 3200 8430 3220 8540
rect 3330 8430 3350 8540
rect 3200 7150 3350 8430
rect 5980 8290 6060 8300
rect 6440 8290 6520 8300
rect 5980 8230 5990 8290
rect 6050 8230 6450 8290
rect 6510 8230 6520 8290
rect 5980 8220 6060 8230
rect 6440 8220 6520 8230
rect 3200 7080 3480 7150
rect 3200 6950 3270 7080
rect 3420 6950 3480 7080
rect 3200 6910 3480 6950
rect 3330 6670 3480 6910
rect 4190 4030 4290 4040
rect 4190 3950 4200 4030
rect 4280 4020 4290 4030
rect 4430 4030 4530 4040
rect 4430 4020 4440 4030
rect 4280 3960 4440 4020
rect 4280 3950 4290 3960
rect 4190 3940 4290 3950
rect 4430 3950 4440 3960
rect 4520 3950 4530 4030
rect 4430 3940 4530 3950
<< via2 >>
rect 4320 12420 4400 12500
rect 6450 8230 6510 8290
rect 3270 6950 3420 7080
rect 4200 3950 4280 4030
<< metal3 >>
rect 340 12500 440 12510
rect 340 12420 350 12500
rect 430 12490 440 12500
rect 4310 12500 4410 12510
rect 4310 12490 4320 12500
rect 430 12430 4320 12490
rect 430 12420 440 12430
rect 340 12410 440 12420
rect 4310 12420 4320 12430
rect 4400 12420 4410 12500
rect 4310 12410 4410 12420
rect 7190 8300 7340 8310
rect 6440 8290 6520 8300
rect 7190 8290 7220 8300
rect 6440 8230 6450 8290
rect 6510 8230 7220 8290
rect 6440 8220 6520 8230
rect 7190 8220 7220 8230
rect 7310 8220 7340 8300
rect 7190 8210 7340 8220
rect 3200 7150 3350 7400
rect 3200 7080 3480 7150
rect 3200 6950 3270 7080
rect 3420 6950 3480 7080
rect 3200 6910 3480 6950
rect 3330 3690 3480 6910
rect 4020 4030 4120 4040
rect 4020 3950 4030 4030
rect 4110 4020 4120 4030
rect 4190 4030 4290 4040
rect 4190 4020 4200 4030
rect 4110 3960 4200 4020
rect 4110 3950 4120 3960
rect 4020 3940 4120 3950
rect 4190 3950 4200 3960
rect 4280 3950 4290 4030
rect 4190 3940 4290 3950
rect 3330 3580 3350 3690
rect 3460 3580 3480 3690
rect 3330 3570 3480 3580
<< via3 >>
rect 350 12420 430 12500
rect 7220 8220 7310 8300
rect 4030 3950 4110 4030
rect 3350 3580 3460 3690
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 18500 600 44152
rect 200 18420 340 18500
rect 420 18420 600 18500
rect 200 12500 600 18420
rect 200 12420 350 12500
rect 430 12420 600 12500
rect 200 1000 600 12420
rect 800 4020 1200 44152
rect 7190 8300 7340 8310
rect 7190 8220 7220 8300
rect 7310 8220 7340 8300
rect 4020 4030 4120 4040
rect 4020 4020 4030 4030
rect 800 3960 4030 4020
rect 800 1000 1200 3960
rect 4020 3950 4030 3960
rect 4110 3950 4120 4030
rect 4020 3940 4120 3950
rect 3330 3690 3480 3710
rect 3330 3580 3350 3690
rect 3460 3580 3480 3690
rect 3330 200 3480 3580
rect 7190 200 7340 8220
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
use sky130_fd_pr__res_high_po_0p35_EB26MW  sky130_fd_pr__res_high_po_0p35_EB26MW_1 /foss/designs
timestamp 1739978212
transform 1 0 3547 0 1 9453
box -35 -623 35 623
use sky130_fd_pr__res_xhigh_po_0p35_JEQFFF  sky130_fd_pr__res_xhigh_po_0p35_JEQFFF_1 /foss/designs
timestamp 1739978212
transform 1 0 4257 0 1 13837
box -35 -5647 35 5647
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 340 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1190 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
rlabel metal1 5442 12430 5462 12490 7 VDD
port 3 w
rlabel viali 5562 8240 5602 8280 3 Vout
port 2 e
rlabel metal1 5422 3960 5442 4020 7 GND
port 4 w
<< properties >>
string (UNNAMED) gencell
string FIXED_BBOX 0 0 32200 45152
<< end >>
