* NGSPICE file created from tt_um_alexandercoabad_mixedsignal.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_TEWFY7 a_208_n400# a_366_n400# a_108_n488# a_50_n400#
+ a_n208_n488# a_266_n488# a_n366_n488# a_n108_n400# a_n266_n400# a_n50_n488# a_n526_n574#
+ a_n424_n400#
X0 a_n266_n400# a_n366_n488# a_n424_n400# a_n526_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_366_n400# a_266_n488# a_208_n400# a_n526_n574# sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2 a_50_n400# a_n50_n488# a_n108_n400# a_n526_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n108_n400# a_n208_n488# a_n266_n400# a_n526_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X4 a_208_n400# a_108_n488# a_50_n400# a_n526_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_X45PJH a_n208_n497# a_266_n497# a_208_n400# a_n366_n497#
+ a_366_n400# a_n50_n497# a_50_n400# w_n562_n619# a_n108_n400# a_n266_n400# a_n424_n400#
+ a_108_n497#
X0 a_n266_n400# a_n366_n497# a_n424_n400# w_n562_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_366_n400# a_266_n497# a_208_n400# w_n562_n619# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2 a_50_n400# a_n50_n497# a_n108_n400# w_n562_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n108_n400# a_n208_n497# a_n266_n400# w_n562_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X4 a_208_n400# a_108_n497# a_50_n400# w_n562_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt Inverter_base m1_330_n303# li_73_1291# m1_260_n192# VSUBS
Xsky130_fd_pr__nfet_01v8_TEWFY7_0 VSUBS m1_330_n303# m1_260_n192# m1_330_n303# m1_260_n192#
+ m1_260_n192# m1_260_n192# VSUBS m1_330_n303# m1_260_n192# VSUBS VSUBS sky130_fd_pr__nfet_01v8_TEWFY7
Xsky130_fd_pr__pfet_01v8_X45PJH_0 m1_260_n192# m1_260_n192# li_73_1291# m1_260_n192#
+ m1_330_n303# m1_260_n192# m1_330_n303# li_73_1291# li_73_1291# m1_330_n303# li_73_1291#
+ m1_260_n192# sky130_fd_pr__pfet_01v8_X45PJH
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_PZF9TG a_n573_n1276# a_n573_844# a_n703_n1406#
X0 a_n573_844# a_n573_n1276# a_n703_n1406# sky130_fd_pr__res_xhigh_po_5p73 l=8.6
.ends

.subckt x300k_res sky130_fd_pr__res_xhigh_po_5p73_PZF9TG_29/a_n573_n1276# sky130_fd_pr__res_xhigh_po_5p73_PZF9TG_11/a_n573_n1276#
+ VSUBS
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_0 m1_5001_39611# m1_5001_42495# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_1 m1_5001_36727# m1_5001_39611# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_2 m1_6479_39611# m1_6479_42495# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_3 m1_7957_39611# m1_7957_42495# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_4 m1_9435_39611# m1_9435_42495# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_90 m1_5001_54031# m1_5001_56915# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_5 m1_6479_36727# m1_6479_39611# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_80 m1_12391_48263# m1_12391_51147# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_91 m1_6479_54031# m1_5001_56915# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_6 m1_7957_36727# m1_7957_39611# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_70 m1_18303_45379# m1_18303_48263# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_81 m1_13869_48263# m1_13869_51147# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_92 m1_7957_54031# m1_7957_56915# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_7 m1_9435_36727# m1_9435_39611# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_82 m1_6479_45379# m1_6479_48263# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_71 m1_18303_48263# m1_18303_51147# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_60 m1_18303_51147# m1_18303_54031# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_93 m1_9435_54031# m1_7957_56915# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_8 m1_10913_39611# m1_10913_42495# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_50 m1_5001_42495# m1_5001_45379# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_83 m1_7957_45379# m1_7957_48263# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_72 m1_15347_45379# m1_15347_48263# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_61 m1_15347_51147# m1_15347_54031# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_94 m1_10913_54031# m1_10913_56915# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_40 m1_13869_33843# m1_13869_36727# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_9 m1_12391_39611# m1_12391_42495# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_51 m1_6479_42495# m1_6479_45379# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_84 m1_9435_45379# m1_9435_48263# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_73 m1_16825_45379# m1_16825_48263# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_62 m1_16825_51147# m1_16825_54031# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_95 m1_12391_54031# m1_10913_56915# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_96 m1_13869_54031# m1_13869_56915# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_41 m1_10913_30959# m1_10913_33843# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_30 m1_5001_33843# m1_5001_36727# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_52 m1_7957_42495# m1_7957_45379# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_85 m1_6479_48263# m1_6479_51147# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_74 m1_15347_48263# m1_15347_51147# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_63 m1_10913_51147# m1_10913_54031# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_97 m1_15347_54031# m1_13869_56915# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_31 m1_5001_30959# m1_5001_33843# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_20 m1_12391_28839# m1_12391_30959# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_42 m1_12391_30959# m1_12391_33843# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_53 m1_9435_42495# m1_9435_45379# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_86 m1_7957_48263# m1_7957_51147# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_75 m1_16825_48263# m1_16825_51147# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_64 m1_12391_51147# m1_12391_54031# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_98 m1_16825_54031# m1_16825_56915# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_21 m1_9435_28839# m1_10913_30959# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_43 m1_13869_30959# m1_13869_33843# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_32 m1_6479_33843# m1_6479_36727# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_10 m1_13869_39611# m1_13869_42495# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_54 m1_10913_42495# m1_10913_45379# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_76 m1_10913_45379# m1_10913_48263# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_87 m1_9435_48263# m1_9435_51147# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_65 m1_13869_51147# m1_13869_54031# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_99 m1_18303_54031# m1_16825_56915# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_11 sky130_fd_pr__res_xhigh_po_5p73_PZF9TG_11/a_n573_n1276#
+ m1_18303_30959# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_33 m1_7957_33843# m1_7957_36727# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_44 m1_15347_33843# m1_15347_36727# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_22 m1_15347_36727# m1_15347_39611# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_55 m1_12391_42495# m1_12391_45379# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_88 m1_5001_45379# m1_5001_48263# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_77 m1_12391_45379# m1_12391_48263# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_66 m1_6479_51147# m1_6479_54031# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_34 m1_9435_33843# m1_9435_36727# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_45 m1_16825_33843# m1_16825_36727# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_12 m1_10913_36727# m1_10913_39611# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_23 m1_16825_36727# m1_16825_39611# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_56 m1_13869_42495# m1_13869_45379# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_78 m1_13869_45379# m1_13869_48263# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_89 m1_5001_48263# m1_5001_51147# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_67 m1_7957_51147# m1_7957_54031# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_35 m1_6479_30959# m1_6479_33843# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_46 m1_15347_30959# m1_15347_33843# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_13 m1_12391_36727# m1_12391_39611# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_24 m1_18303_39611# m1_18303_42495# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_57 m1_15347_42495# m1_15347_45379# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_79 m1_10913_48263# m1_10913_51147# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_68 m1_9435_51147# m1_9435_54031# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_14 m1_15347_28839# m1_16825_30959# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_36 m1_7957_30959# m1_7957_33843# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_25 m1_9435_28839# m1_9435_30959# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_47 m1_16825_30959# m1_16825_33843# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_58 m1_16825_42495# m1_16825_45379# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_69 m1_5001_51147# m1_5001_54031# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_26 m1_6479_28839# m1_7957_30959# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_37 m1_9435_30959# m1_9435_33843# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_15 m1_15347_28839# m1_15347_30959# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_48 m1_18303_33843# m1_18303_36727# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_59 m1_18303_42495# m1_18303_45379# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_27 m1_6479_28839# m1_6479_30959# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_49 m1_18303_30959# m1_18303_33843# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_38 m1_10913_33843# m1_10913_36727# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_16 m1_13869_36727# m1_13869_39611# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_39 m1_12391_33843# m1_12391_36727# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_28 m1_18303_36727# m1_18303_39611# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_17 m1_15347_39611# m1_15347_42495# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_29 sky130_fd_pr__res_xhigh_po_5p73_PZF9TG_29/a_n573_n1276#
+ m1_5001_30959# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_18 m1_16825_39611# m1_16825_42495# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_19 m1_12391_28839# m1_13869_30959# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
.ends

.subckt x3k_res XR3/a_n573_844# XR3/a_n573_n1276# VSUBS
XXR3 XR3/a_n573_n1276# XR3/a_n573_844# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
.ends

.subckt sky130_fd_pr__nfet_01v8_JZTGL9 a_n260_n274# a_100_n100# a_n158_n100# a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n260_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_U6BDKB w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt Inverter Vin Vout VDD GND
Xsky130_fd_pr__nfet_01v8_JZTGL9_0 GND Vout GND Vin sky130_fd_pr__nfet_01v8_JZTGL9
Xsky130_fd_pr__pfet_01v8_U6BDKB_0 VDD Vin Vout VDD sky130_fd_pr__pfet_01v8_U6BDKB
.ends

.subckt x4-to-1_analog_MUX I1 I2 I3 I4 S1 S2 OUT VDD GND
Xsky130_fd_pr__nfet_01v8_JZTGL9_0 GND m1_278_n644# I1 Inverter_1/Vout sky130_fd_pr__nfet_01v8_JZTGL9
Xsky130_fd_pr__nfet_01v8_JZTGL9_1 GND I4 m1_278_n2780# S1 sky130_fd_pr__nfet_01v8_JZTGL9
Xsky130_fd_pr__nfet_01v8_JZTGL9_2 GND m1_278_n2780# I2 Inverter_1/Vout sky130_fd_pr__nfet_01v8_JZTGL9
Xsky130_fd_pr__nfet_01v8_JZTGL9_3 GND OUT m1_278_n644# S2bar sky130_fd_pr__nfet_01v8_JZTGL9
Xsky130_fd_pr__nfet_01v8_JZTGL9_4 GND I3 m1_278_n644# S1 sky130_fd_pr__nfet_01v8_JZTGL9
Xsky130_fd_pr__nfet_01v8_JZTGL9_5 GND OUT m1_278_n2780# S2 sky130_fd_pr__nfet_01v8_JZTGL9
Xsky130_fd_pr__pfet_01v8_U6BDKB_0 VDD S2 OUT m1_278_n644# sky130_fd_pr__pfet_01v8_U6BDKB
Xsky130_fd_pr__pfet_01v8_U6BDKB_1 VDD Inverter_1/Vout I4 m1_278_n2780# sky130_fd_pr__pfet_01v8_U6BDKB
Xsky130_fd_pr__pfet_01v8_U6BDKB_2 VDD S1 m1_278_n2780# I2 sky130_fd_pr__pfet_01v8_U6BDKB
Xsky130_fd_pr__pfet_01v8_U6BDKB_3 VDD S1 m1_278_n644# I1 sky130_fd_pr__pfet_01v8_U6BDKB
Xsky130_fd_pr__pfet_01v8_U6BDKB_4 VDD Inverter_1/Vout I3 m1_278_n644# sky130_fd_pr__pfet_01v8_U6BDKB
Xsky130_fd_pr__pfet_01v8_U6BDKB_5 VDD S2bar OUT m1_278_n2780# sky130_fd_pr__pfet_01v8_U6BDKB
XInverter_1 S1 Inverter_1/Vout VDD GND Inverter
XInverter_0 S2 S2bar VDD GND Inverter
.ends

.subckt x30k_res sky130_fd_pr__res_xhigh_po_5p73_PZF9TG_0/a_n573_n1276# sky130_fd_pr__res_xhigh_po_5p73_PZF9TG_3/a_n573_n1276#
+ VSUBS
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_0 sky130_fd_pr__res_xhigh_po_5p73_PZF9TG_0/a_n573_n1276#
+ m1_11905_2235# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_1 m1_10427_115# m1_11905_2235# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_2 m1_1559_115# m1_81_2235# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_3 sky130_fd_pr__res_xhigh_po_5p73_PZF9TG_3/a_n573_n1276#
+ m1_81_2235# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_4 m1_7471_115# m1_8949_2235# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_5 m1_10427_115# m1_8949_2235# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_7 m1_7471_115# m1_5993_2235# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_6 m1_4515_115# m1_5993_2235# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_8 m1_1559_115# m1_3037_2235# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
Xsky130_fd_pr__res_xhigh_po_5p73_PZF9TG_9 m1_4515_115# m1_3037_2235# VSUBS sky130_fd_pr__res_xhigh_po_5p73_PZF9TG
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_UP82F9 a_n573_n703# a_n703_n833# a_n573_271#
X0 a_n573_271# a_n573_n703# a_n703_n833# sky130_fd_pr__res_xhigh_po_5p73 l=2.87
.ends

.subckt x100k_res sky130_fd_pr__res_xhigh_po_5p73_UP82F9_7/a_n573_n703# sky130_fd_pr__res_xhigh_po_5p73_UP82F9_0/a_n573_n703#
+ VSUBS
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_8 m1_10425_119# VSUBS m1_10425_1093# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_9 m1_7469_119# VSUBS m1_8947_1093# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_90 m1_79_14997# VSUBS m1_79_16735# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_80 m1_1557_13259# VSUBS m1_1557_14997# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_91 m1_1557_14997# VSUBS m1_79_16735# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_70 m1_13381_9783# VSUBS m1_13381_11521# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_81 m1_79_13259# VSUBS m1_79_14997# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_92 m1_3035_14997# VSUBS m1_3035_16735# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_71 m1_11903_9783# VSUBS m1_11903_11521# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_60 m1_13381_11521# VSUBS m1_13381_13259# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_82 m1_4513_13259# VSUBS m1_4513_14997# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_93 m1_4513_14997# VSUBS m1_3035_16735# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_50 m1_7469_6307# VSUBS m1_7469_8045# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_72 m1_10425_9783# VSUBS m1_10425_11521# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_61 m1_8947_11521# VSUBS m1_8947_13259# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_83 m1_3035_13259# VSUBS m1_3035_14997# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_94 m1_5991_14997# VSUBS m1_5991_16735# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_51 m1_5991_6307# VSUBS m1_5991_8045# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_40 m1_79_8045# VSUBS m1_79_9783# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_73 m1_8947_9783# VSUBS m1_8947_11521# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_62 m1_10425_11521# VSUBS m1_10425_13259# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_84 m1_7469_13259# VSUBS m1_7469_14997# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_95 m1_7469_14997# VSUBS m1_5991_16735# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_96 m1_8947_14997# VSUBS m1_8947_16735# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_30 m1_13381_4569# VSUBS m1_13381_6307# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_41 m1_1557_8045# VSUBS m1_1557_9783# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_52 m1_8947_8045# VSUBS m1_8947_9783# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_74 m1_7469_9783# VSUBS m1_7469_11521# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_63 m1_11903_11521# VSUBS m1_11903_13259# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_85 m1_5991_13259# VSUBS m1_5991_14997# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_97 m1_10425_14997# VSUBS m1_8947_16735# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_20 m1_1557_2831# VSUBS m1_1557_4569# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_31 m1_8947_4569# VSUBS m1_8947_6307# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_42 m1_1557_6307# VSUBS m1_1557_8045# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_53 m1_10425_8045# VSUBS m1_10425_9783# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_75 m1_5991_9783# VSUBS m1_5991_11521# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_64 m1_5991_11521# VSUBS m1_5991_13259# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_86 m1_11903_13259# VSUBS m1_11903_14997# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_98 m1_11903_14997# VSUBS m1_11903_16735# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_10 m1_13381_1093# VSUBS m1_13381_2831# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_21 m1_79_2831# VSUBS m1_79_4569# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_32 m1_10425_4569# VSUBS m1_10425_6307# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_43 m1_79_6307# VSUBS m1_79_8045# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_54 m1_11903_8045# VSUBS m1_11903_9783# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_76 m1_4513_9783# VSUBS m1_4513_11521# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_65 m1_7469_11521# VSUBS m1_7469_13259# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_87 m1_10425_13259# VSUBS m1_10425_14997# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_99 m1_13381_14997# VSUBS m1_11903_16735# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_11 m1_11903_1093# VSUBS m1_11903_2831# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_22 m1_4513_2831# VSUBS m1_4513_4569# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_33 m1_11903_4569# VSUBS m1_11903_6307# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_55 m1_11903_6307# VSUBS m1_11903_8045# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_44 m1_3035_8045# VSUBS m1_3035_9783# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_77 m1_3035_9783# VSUBS m1_3035_11521# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_66 m1_3035_11521# VSUBS m1_3035_13259# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_88 m1_8947_13259# VSUBS m1_8947_14997# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_12 m1_10425_1093# VSUBS m1_10425_2831# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_23 m1_3035_2831# VSUBS m1_3035_4569# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_34 m1_5991_4569# VSUBS m1_5991_6307# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_56 m1_10425_6307# VSUBS m1_10425_8045# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_45 m1_4513_8045# VSUBS m1_4513_9783# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_78 m1_1557_9783# VSUBS m1_1557_11521# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_67 m1_4513_11521# VSUBS m1_4513_13259# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_89 m1_13381_13259# VSUBS m1_13381_14997# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_13 m1_8947_1093# VSUBS m1_8947_2831# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_24 m1_7469_2831# VSUBS m1_7469_4569# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_35 m1_7469_4569# VSUBS m1_7469_6307# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_46 m1_4513_6307# VSUBS m1_4513_8045# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_57 m1_8947_6307# VSUBS m1_8947_8045# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_79 m1_79_9783# VSUBS m1_79_11521# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_68 m1_79_11521# VSUBS m1_79_13259# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_14 m1_7469_1093# VSUBS m1_7469_2831# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_0 sky130_fd_pr__res_xhigh_po_5p73_UP82F9_0/a_n573_n703#
+ VSUBS m1_13381_1093# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_25 m1_5991_2831# VSUBS m1_5991_4569# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_36 m1_3035_4569# VSUBS m1_3035_6307# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_47 m1_3035_6307# VSUBS m1_3035_8045# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_58 m1_13381_8045# VSUBS m1_13381_9783# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_69 m1_1557_11521# VSUBS m1_1557_13259# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_1 m1_10425_119# VSUBS m1_11903_1093# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_15 m1_5991_1093# VSUBS m1_5991_2831# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_26 m1_11903_2831# VSUBS m1_11903_4569# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_37 m1_4513_4569# VSUBS m1_4513_6307# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_59 m1_13381_6307# VSUBS m1_13381_8045# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_48 m1_5991_8045# VSUBS m1_5991_9783# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_16 m1_4513_1093# VSUBS m1_4513_2831# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_2 m1_7469_119# VSUBS m1_7469_1093# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_27 m1_10425_2831# VSUBS m1_10425_4569# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_38 m1_79_4569# VSUBS m1_79_6307# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_49 m1_7469_8045# VSUBS m1_7469_9783# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_17 m1_3035_1093# VSUBS m1_3035_2831# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_3 m1_4513_119# VSUBS m1_5991_1093# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_28 m1_8947_2831# VSUBS m1_8947_4569# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_39 m1_1557_4569# VSUBS m1_1557_6307# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_18 m1_1557_1093# VSUBS m1_1557_2831# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_4 m1_1557_119# VSUBS m1_3035_1093# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_29 m1_13381_2831# VSUBS m1_13381_4569# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_19 m1_79_1093# VSUBS m1_79_2831# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_5 m1_4513_119# VSUBS m1_4513_1093# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_6 m1_1557_119# VSUBS m1_1557_1093# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
Xsky130_fd_pr__res_xhigh_po_5p73_UP82F9_7 sky130_fd_pr__res_xhigh_po_5p73_UP82F9_7/a_n573_n703#
+ VSUBS m1_79_1093# sky130_fd_pr__res_xhigh_po_5p73_UP82F9
.ends

.subckt tt_um_alexandercoabad_mixedsignal clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4]
+ ua[5] ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6]
+ ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VDPWR VGND
XInverter_base_0 ua[0] VDPWR mux_in VGND Inverter_base
X300k_res_1 ua[0] mux_in VGND x300k_res
X3k_res_0 3k_res_0/XR3/a_n573_844# mux_in VGND x3k_res
X3k_res_1 4-to-1_analog_MUX_0/I3 ua[0] VGND x3k_res
X4-to-1_analog_MUX_0 4-to-1_analog_MUX_0/I1 4-to-1_analog_MUX_0/I2 4-to-1_analog_MUX_0/I3
+ 4-to-1_analog_MUX_0/I4 4-to-1_analog_MUX_0/S1 4-to-1_analog_MUX_0/S2 mux_in VDPWR
+ VGND x4-to-1_analog_MUX
X30k_res_0 ua[0] 4-to-1_analog_MUX_0/I2 VGND x30k_res
X100k_res_1 4-to-1_analog_MUX_0/I4 ua[0] VGND x100k_res
.ends

