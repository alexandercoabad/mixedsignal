magic
tech sky130A
magscale 1 2
timestamp 1757858607
<< nwell >>
rect -562 -619 562 619
<< pmos >>
rect -366 -400 -266 400
rect -208 -400 -108 400
rect -50 -400 50 400
rect 108 -400 208 400
rect 266 -400 366 400
<< pdiff >>
rect -424 388 -366 400
rect -424 -388 -412 388
rect -378 -388 -366 388
rect -424 -400 -366 -388
rect -266 388 -208 400
rect -266 -388 -254 388
rect -220 -388 -208 388
rect -266 -400 -208 -388
rect -108 388 -50 400
rect -108 -388 -96 388
rect -62 -388 -50 388
rect -108 -400 -50 -388
rect 50 388 108 400
rect 50 -388 62 388
rect 96 -388 108 388
rect 50 -400 108 -388
rect 208 388 266 400
rect 208 -388 220 388
rect 254 -388 266 388
rect 208 -400 266 -388
rect 366 388 424 400
rect 366 -388 378 388
rect 412 -388 424 388
rect 366 -400 424 -388
<< pdiffc >>
rect -412 -388 -378 388
rect -254 -388 -220 388
rect -96 -388 -62 388
rect 62 -388 96 388
rect 220 -388 254 388
rect 378 -388 412 388
<< nsubdiff >>
rect -526 549 -430 583
rect 430 549 526 583
rect -526 487 -492 549
rect 492 487 526 549
rect -526 -549 -492 -487
rect 492 -549 526 -487
rect -526 -583 -430 -549
rect 430 -583 526 -549
<< nsubdiffcont >>
rect -430 549 430 583
rect -526 -487 -492 487
rect 492 -487 526 487
rect -430 -583 430 -549
<< poly >>
rect -366 400 -266 497
rect -208 400 -108 497
rect -50 400 50 497
rect 108 400 208 497
rect 266 400 366 497
rect -366 -447 -266 -400
rect -366 -481 -350 -447
rect -282 -481 -266 -447
rect -366 -497 -266 -481
rect -208 -447 -108 -400
rect -208 -481 -192 -447
rect -124 -481 -108 -447
rect -208 -497 -108 -481
rect -50 -447 50 -400
rect -50 -481 -34 -447
rect 34 -481 50 -447
rect -50 -497 50 -481
rect 108 -447 208 -400
rect 108 -481 124 -447
rect 192 -481 208 -447
rect 108 -497 208 -481
rect 266 -447 366 -400
rect 266 -481 282 -447
rect 350 -481 366 -447
rect 266 -497 366 -481
<< polycont >>
rect -350 -481 -282 -447
rect -192 -481 -124 -447
rect -34 -481 34 -447
rect 124 -481 192 -447
rect 282 -481 350 -447
<< locali >>
rect -526 549 -430 583
rect 430 549 526 583
rect -526 487 -492 549
rect 492 487 526 549
rect -412 388 -378 404
rect -412 -404 -378 -388
rect -254 388 -220 404
rect -254 -404 -220 -388
rect -96 388 -62 404
rect -96 -404 -62 -388
rect 62 388 96 404
rect 62 -404 96 -388
rect 220 388 254 404
rect 220 -404 254 -388
rect 378 388 412 404
rect 378 -404 412 -388
rect -366 -481 -350 -447
rect -282 -481 -266 -447
rect -208 -481 -192 -447
rect -124 -481 -108 -447
rect -50 -481 -34 -447
rect 34 -481 50 -447
rect 108 -481 124 -447
rect 192 -481 208 -447
rect 266 -481 282 -447
rect 350 -481 366 -447
rect -526 -549 -492 -487
rect 492 -549 526 -487
rect -526 -583 -430 -549
rect 430 -583 526 -549
<< viali >>
rect -412 -388 -378 388
rect -254 -388 -220 388
rect -96 -388 -62 388
rect 62 -388 96 388
rect 220 -388 254 388
rect 378 -388 412 388
rect -350 -481 -282 -447
rect -192 -481 -124 -447
rect -34 -481 34 -447
rect 124 -481 192 -447
rect 282 -481 350 -447
<< metal1 >>
rect -418 388 -372 400
rect -418 -388 -412 388
rect -378 -388 -372 388
rect -418 -400 -372 -388
rect -260 388 -214 400
rect -260 -388 -254 388
rect -220 -388 -214 388
rect -260 -400 -214 -388
rect -102 388 -56 400
rect -102 -388 -96 388
rect -62 -388 -56 388
rect -102 -400 -56 -388
rect 56 388 102 400
rect 56 -388 62 388
rect 96 -388 102 388
rect 56 -400 102 -388
rect 214 388 260 400
rect 214 -388 220 388
rect 254 -388 260 388
rect 214 -400 260 -388
rect 372 388 418 400
rect 372 -388 378 388
rect 412 -388 418 388
rect 372 -400 418 -388
rect -362 -447 -270 -441
rect -362 -481 -350 -447
rect -282 -481 -270 -447
rect -362 -487 -270 -481
rect -204 -447 -112 -441
rect -204 -481 -192 -447
rect -124 -481 -112 -447
rect -204 -487 -112 -481
rect -46 -447 46 -441
rect -46 -481 -34 -447
rect 34 -481 46 -447
rect -46 -487 46 -481
rect 112 -447 204 -441
rect 112 -481 124 -447
rect 192 -481 204 -447
rect 112 -487 204 -481
rect 270 -447 362 -441
rect 270 -481 282 -447
rect 350 -481 362 -447
rect 270 -487 362 -481
<< properties >>
string FIXED_BBOX -509 -566 509 566
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4 l 0.5 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__pfet_01v8_X45PJH parameters
<< end >>
