magic
tech sky130A
magscale 1 2
timestamp 1740568496
<< nwell >>
rect 27942 8290 28644 12510
<< nmos >>
rect 28282 4050 28382 8050
<< pmos >>
rect 28282 8400 28382 12400
<< ndiff >>
rect 28062 8020 28282 8050
rect 28062 4080 28152 8020
rect 28192 4080 28282 8020
rect 28062 4050 28282 4080
rect 28382 8020 28602 8050
rect 28382 4080 28472 8020
rect 28512 4080 28602 8020
rect 28382 4050 28602 4080
<< pdiff >>
rect 28062 12370 28282 12400
rect 28062 8430 28152 12370
rect 28192 8430 28282 12370
rect 28062 8400 28282 8430
rect 28382 12370 28602 12400
rect 28382 8430 28472 12370
rect 28512 8430 28602 12370
rect 28382 8400 28602 8430
<< ndiffc >>
rect 28152 4080 28192 8020
rect 28472 4080 28512 8020
<< pdiffc >>
rect 28152 8430 28192 12370
rect 28472 8430 28512 12370
<< psubdiff >>
rect 27982 8020 28062 8050
rect 27982 4080 28002 8020
rect 28042 4080 28062 8020
rect 27982 4050 28062 4080
<< nsubdiff >>
rect 27982 12370 28062 12400
rect 27982 8430 28002 12370
rect 28042 8430 28062 12370
rect 27982 8400 28062 8430
<< psubdiffcont >>
rect 28002 4080 28042 8020
<< nsubdiffcont >>
rect 28002 8430 28042 12370
<< poly >>
rect 28282 12400 28382 12500
rect 28282 8290 28382 8400
rect 28202 8280 28382 8290
rect 28202 8240 28222 8280
rect 28262 8240 28382 8280
rect 28202 8230 28382 8240
rect 28282 8050 28382 8230
rect 28282 3950 28382 4050
<< polycont >>
rect 28222 8240 28262 8280
<< locali >>
rect 27982 12390 28022 12440
rect 27982 12370 28272 12390
rect 27982 8430 28002 12370
rect 28042 8430 28152 12370
rect 28192 8430 28272 12370
rect 27982 8410 28272 8430
rect 28392 12370 28602 12390
rect 28392 8430 28472 12370
rect 28512 8430 28602 12370
rect 28392 8290 28602 8430
rect 27922 8280 28282 8290
rect 27922 8240 27942 8280
rect 27982 8240 28222 8280
rect 28262 8240 28282 8280
rect 27922 8230 28282 8240
rect 28392 8280 28802 8290
rect 28392 8240 28740 8280
rect 28790 8240 28802 8280
rect 28392 8230 28802 8240
rect 27982 8020 28272 8040
rect 27982 4080 28002 8020
rect 28042 4080 28152 8020
rect 28192 4080 28272 8020
rect 27982 4060 28272 4080
rect 28392 8020 28602 8230
rect 28392 4080 28472 8020
rect 28512 4080 28602 8020
rect 28392 4060 28602 4080
rect 27982 4010 28022 4060
<< viali >>
rect 27980 12440 28022 12480
rect 27942 8240 27982 8280
rect 28740 8240 28790 8280
rect 27982 3970 28022 4010
<< metal1 >>
rect 27432 19130 28792 19200
rect 27680 12430 27700 12490
rect 27760 12480 28610 12490
rect 27760 12440 27980 12480
rect 28022 12440 28610 12480
rect 27760 12430 28610 12440
rect 26380 9870 26760 9940
rect 26380 8540 26530 9870
rect 26380 8430 26400 8540
rect 26510 8430 26530 8540
rect 26692 8290 26762 8890
rect 28722 8290 28792 19130
rect 29160 8290 29240 8300
rect 26692 8280 28002 8290
rect 26692 8240 27942 8280
rect 27982 8240 28002 8280
rect 26692 8230 28002 8240
rect 28720 8280 29170 8290
rect 28720 8240 28740 8280
rect 28790 8240 29170 8280
rect 28720 8230 29170 8240
rect 29230 8230 29240 8290
rect 29160 8220 29240 8230
rect 27610 4030 27710 4040
rect 27610 3950 27620 4030
rect 27700 4020 27710 4030
rect 27700 4010 28590 4020
rect 27700 3970 27982 4010
rect 28022 3970 28590 4010
rect 27700 3960 28590 3970
rect 27700 3950 27710 3960
rect 27610 3940 27710 3950
<< via1 >>
rect 27700 12430 27760 12490
rect 26400 8430 26510 8540
rect 29170 8230 29230 8290
rect 27620 3950 27700 4030
<< metal2 >>
rect 27490 12500 27590 12510
rect 27490 12420 27500 12500
rect 27580 12490 27590 12500
rect 27580 12430 27700 12490
rect 27760 12430 27770 12490
rect 27580 12420 27590 12430
rect 27490 12410 27590 12420
rect 26380 8540 26530 8550
rect 26380 8430 26400 8540
rect 26510 8430 26530 8540
rect 26380 7150 26530 8430
rect 29160 8290 29240 8300
rect 29620 8290 29700 8300
rect 29160 8230 29170 8290
rect 29230 8230 29630 8290
rect 29690 8230 29700 8290
rect 29160 8220 29240 8230
rect 29620 8220 29700 8230
rect 26380 7080 26660 7150
rect 26380 6950 26450 7080
rect 26600 6950 26660 7080
rect 26380 6910 26660 6950
rect 26510 6670 26660 6910
rect 27370 4030 27470 4040
rect 27370 3950 27380 4030
rect 27460 4020 27470 4030
rect 27610 4030 27710 4040
rect 27610 4020 27620 4030
rect 27460 3960 27620 4020
rect 27460 3950 27470 3960
rect 27370 3940 27470 3950
rect 27610 3950 27620 3960
rect 27700 3950 27710 4030
rect 27610 3940 27710 3950
<< via2 >>
rect 27500 12420 27580 12500
rect 29630 8230 29690 8290
rect 26450 6950 26600 7080
rect 27380 3950 27460 4030
<< metal3 >>
rect 320 12510 440 12520
rect 320 12490 330 12510
rect 310 12430 330 12490
rect 320 12410 330 12430
rect 430 12490 440 12510
rect 27490 12500 27590 12510
rect 27490 12490 27500 12500
rect 430 12430 27500 12490
rect 430 12410 440 12430
rect 27490 12420 27500 12430
rect 27580 12420 27590 12500
rect 27490 12410 27590 12420
rect 320 12400 440 12410
rect 30370 8300 30520 8310
rect 29620 8290 29700 8300
rect 30370 8290 30400 8300
rect 29620 8230 29630 8290
rect 29690 8230 30400 8290
rect 29620 8220 29700 8230
rect 30370 8220 30400 8230
rect 30490 8220 30520 8300
rect 30370 8210 30520 8220
rect 26380 7150 26530 7400
rect 26380 7080 26660 7150
rect 26380 6950 26450 7080
rect 26600 6950 26660 7080
rect 26380 6910 26660 6950
rect 26510 3690 26660 6910
rect 27200 4030 27300 4040
rect 27200 3950 27210 4030
rect 27290 4020 27300 4030
rect 27370 4030 27470 4040
rect 27370 4020 27380 4030
rect 27290 3960 27380 4020
rect 27290 3950 27300 3960
rect 27200 3940 27300 3950
rect 27370 3950 27380 3960
rect 27460 3950 27470 4030
rect 27370 3940 27470 3950
rect 26510 3580 26530 3690
rect 26640 3580 26660 3690
rect 26510 3570 26660 3580
<< via3 >>
rect 330 12410 430 12510
rect 30400 8220 30490 8300
rect 27210 3950 27290 4030
rect 26530 3580 26640 3690
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 12510 600 44152
rect 200 12410 330 12510
rect 430 12410 600 12510
rect 200 1000 600 12410
rect 800 4020 1200 44152
rect 30370 8300 30520 8310
rect 30370 8220 30400 8300
rect 30490 8220 30520 8300
rect 27200 4030 27300 4040
rect 27200 4020 27210 4030
rect 800 3960 27210 4020
rect 800 1000 1200 3960
rect 27200 3950 27210 3960
rect 27290 3950 27300 4030
rect 27200 3940 27300 3950
rect 26510 3690 26660 3710
rect 26510 3580 26530 3690
rect 26640 3580 26660 3690
rect 26510 200 26660 3580
rect 30370 200 30520 8220
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
use sky130_fd_pr__res_high_po_0p35_EB26MW  sky130_fd_pr__res_high_po_0p35_EB26MW_1 /foss/designs
timestamp 1739978212
transform 1 0 26727 0 1 9453
box -35 -623 35 623
use sky130_fd_pr__res_xhigh_po_0p35_JEQFFF  sky130_fd_pr__res_xhigh_po_0p35_JEQFFF_1 /foss/designs
timestamp 1739978212
transform 1 0 27437 0 1 13837
box -35 -5647 35 5647
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string (UNNAMED) gencell
string FIXED_BBOX 0 0 32200 45152
<< end >>
