* NGSPICE file created from Inverter.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_JZTGL9 a_n260_n274# a_100_n100# a_n158_n100# a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n260_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_U6BDKB w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt Inverter Vin Vout GND VDD
Xsky130_fd_pr__nfet_01v8_JZTGL9_0 GND Vout GND Vin sky130_fd_pr__nfet_01v8_JZTGL9
Xsky130_fd_pr__pfet_01v8_U6BDKB_0 VDD Vin Vout VDD sky130_fd_pr__pfet_01v8_U6BDKB
.ends

