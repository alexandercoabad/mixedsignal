VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_alexandercoabad_mixedsignal
  CLASS BLOCK ;
  FOREIGN tt_um_alexandercoabad_mixedsignal ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.960000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.000000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.500000 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 6.130 23.690 80.030 110.590 ;
        RECT 80.180 23.705 154.080 167.905 ;
        RECT 10.760 4.980 84.660 19.400 ;
        RECT 90.605 4.255 97.995 18.675 ;
      LAYER nwell ;
        RECT 102.795 16.260 114.635 19.450 ;
      LAYER pwell ;
        RECT 102.795 12.475 114.635 15.575 ;
        RECT 102.795 8.685 114.635 11.785 ;
      LAYER nwell ;
        RECT 102.795 4.810 114.635 8.000 ;
      LAYER pwell ;
        RECT 129.245 2.905 136.635 17.325 ;
      LAYER nwell ;
        RECT 144.420 14.130 150.040 20.320 ;
      LAYER pwell ;
        RECT 144.420 7.345 150.040 13.445 ;
      LAYER li1 ;
        RECT 79.850 167.555 153.900 167.725 ;
        RECT 79.850 153.835 80.530 167.555 ;
        RECT 81.010 164.915 86.740 167.075 ;
        RECT 81.010 154.315 86.740 156.475 ;
        RECT 87.220 153.835 87.390 167.555 ;
        RECT 87.750 153.835 87.920 167.555 ;
        RECT 88.400 164.915 94.130 167.075 ;
        RECT 88.400 154.315 94.130 156.475 ;
        RECT 94.610 153.835 94.780 167.555 ;
        RECT 95.140 153.835 95.310 167.555 ;
        RECT 95.790 164.915 101.520 167.075 ;
        RECT 95.790 154.315 101.520 156.475 ;
        RECT 102.000 153.835 102.170 167.555 ;
        RECT 102.530 153.835 102.700 167.555 ;
        RECT 103.180 164.915 108.910 167.075 ;
        RECT 103.180 154.315 108.910 156.475 ;
        RECT 109.390 153.835 109.560 167.555 ;
        RECT 109.920 153.835 110.090 167.555 ;
        RECT 110.570 164.915 116.300 167.075 ;
        RECT 110.570 154.315 116.300 156.475 ;
        RECT 116.780 153.835 116.950 167.555 ;
        RECT 117.310 153.835 117.480 167.555 ;
        RECT 117.960 164.915 123.690 167.075 ;
        RECT 117.960 154.315 123.690 156.475 ;
        RECT 124.170 153.835 124.340 167.555 ;
        RECT 124.700 153.835 124.870 167.555 ;
        RECT 125.350 164.915 131.080 167.075 ;
        RECT 125.350 154.315 131.080 156.475 ;
        RECT 131.560 153.835 131.730 167.555 ;
        RECT 132.090 153.835 132.260 167.555 ;
        RECT 132.740 164.915 138.470 167.075 ;
        RECT 132.740 154.315 138.470 156.475 ;
        RECT 138.950 153.835 139.120 167.555 ;
        RECT 139.480 153.835 139.650 167.555 ;
        RECT 140.130 164.915 145.860 167.075 ;
        RECT 140.130 154.315 145.860 156.475 ;
        RECT 146.340 153.835 146.510 167.555 ;
        RECT 146.870 153.835 147.040 167.555 ;
        RECT 147.520 164.915 153.250 167.075 ;
        RECT 147.520 154.315 153.250 156.475 ;
        RECT 153.730 153.835 153.900 167.555 ;
        RECT 79.850 153.135 153.900 153.835 ;
        RECT 79.850 139.415 80.530 153.135 ;
        RECT 81.010 150.495 86.740 152.655 ;
        RECT 81.010 139.895 86.740 142.055 ;
        RECT 87.220 139.415 87.390 153.135 ;
        RECT 87.750 139.415 87.920 153.135 ;
        RECT 88.400 150.495 94.130 152.655 ;
        RECT 88.400 139.895 94.130 142.055 ;
        RECT 94.610 139.415 94.780 153.135 ;
        RECT 95.140 139.415 95.310 153.135 ;
        RECT 95.790 150.495 101.520 152.655 ;
        RECT 95.790 139.895 101.520 142.055 ;
        RECT 102.000 139.415 102.170 153.135 ;
        RECT 102.530 139.415 102.700 153.135 ;
        RECT 103.180 150.495 108.910 152.655 ;
        RECT 103.180 139.895 108.910 142.055 ;
        RECT 109.390 139.415 109.560 153.135 ;
        RECT 109.920 139.415 110.090 153.135 ;
        RECT 110.570 150.495 116.300 152.655 ;
        RECT 110.570 139.895 116.300 142.055 ;
        RECT 116.780 139.415 116.950 153.135 ;
        RECT 117.310 139.415 117.480 153.135 ;
        RECT 117.960 150.495 123.690 152.655 ;
        RECT 117.960 139.895 123.690 142.055 ;
        RECT 124.170 139.415 124.340 153.135 ;
        RECT 124.700 139.415 124.870 153.135 ;
        RECT 125.350 150.495 131.080 152.655 ;
        RECT 125.350 139.895 131.080 142.055 ;
        RECT 131.560 139.415 131.730 153.135 ;
        RECT 132.090 139.415 132.260 153.135 ;
        RECT 132.740 150.495 138.470 152.655 ;
        RECT 132.740 139.895 138.470 142.055 ;
        RECT 138.950 139.415 139.120 153.135 ;
        RECT 139.480 139.415 139.650 153.135 ;
        RECT 140.130 150.495 145.860 152.655 ;
        RECT 140.130 139.895 145.860 142.055 ;
        RECT 146.340 139.415 146.510 153.135 ;
        RECT 146.870 139.415 147.040 153.135 ;
        RECT 147.520 150.495 153.250 152.655 ;
        RECT 147.520 139.895 153.250 142.055 ;
        RECT 153.730 139.415 153.900 153.135 ;
        RECT 79.850 138.715 153.900 139.415 ;
        RECT 79.850 124.995 80.530 138.715 ;
        RECT 81.010 136.075 86.740 138.235 ;
        RECT 81.010 125.475 86.740 127.635 ;
        RECT 87.220 124.995 87.390 138.715 ;
        RECT 87.750 124.995 87.920 138.715 ;
        RECT 88.400 136.075 94.130 138.235 ;
        RECT 88.400 125.475 94.130 127.635 ;
        RECT 94.610 124.995 94.780 138.715 ;
        RECT 95.140 124.995 95.310 138.715 ;
        RECT 95.790 136.075 101.520 138.235 ;
        RECT 95.790 125.475 101.520 127.635 ;
        RECT 102.000 124.995 102.170 138.715 ;
        RECT 102.530 124.995 102.700 138.715 ;
        RECT 103.180 136.075 108.910 138.235 ;
        RECT 103.180 125.475 108.910 127.635 ;
        RECT 109.390 124.995 109.560 138.715 ;
        RECT 109.920 124.995 110.090 138.715 ;
        RECT 110.570 136.075 116.300 138.235 ;
        RECT 110.570 125.475 116.300 127.635 ;
        RECT 116.780 124.995 116.950 138.715 ;
        RECT 117.310 124.995 117.480 138.715 ;
        RECT 117.960 136.075 123.690 138.235 ;
        RECT 117.960 125.475 123.690 127.635 ;
        RECT 124.170 124.995 124.340 138.715 ;
        RECT 124.700 124.995 124.870 138.715 ;
        RECT 125.350 136.075 131.080 138.235 ;
        RECT 125.350 125.475 131.080 127.635 ;
        RECT 131.560 124.995 131.730 138.715 ;
        RECT 132.090 124.995 132.260 138.715 ;
        RECT 132.740 136.075 138.470 138.235 ;
        RECT 132.740 125.475 138.470 127.635 ;
        RECT 138.950 124.995 139.120 138.715 ;
        RECT 139.480 124.995 139.650 138.715 ;
        RECT 140.130 136.075 145.860 138.235 ;
        RECT 140.130 125.475 145.860 127.635 ;
        RECT 146.340 124.995 146.510 138.715 ;
        RECT 146.870 124.995 147.040 138.715 ;
        RECT 147.520 136.075 153.250 138.235 ;
        RECT 147.520 125.475 153.250 127.635 ;
        RECT 153.730 124.995 153.900 138.715 ;
        RECT 79.850 124.295 153.900 124.995 ;
        RECT 79.850 110.575 80.530 124.295 ;
        RECT 81.010 121.655 86.740 123.815 ;
        RECT 81.010 111.055 86.740 113.215 ;
        RECT 87.220 110.575 87.390 124.295 ;
        RECT 87.750 110.575 87.920 124.295 ;
        RECT 88.400 121.655 94.130 123.815 ;
        RECT 88.400 111.055 94.130 113.215 ;
        RECT 94.610 110.575 94.780 124.295 ;
        RECT 95.140 110.575 95.310 124.295 ;
        RECT 95.790 121.655 101.520 123.815 ;
        RECT 95.790 111.055 101.520 113.215 ;
        RECT 102.000 110.575 102.170 124.295 ;
        RECT 102.530 110.575 102.700 124.295 ;
        RECT 103.180 121.655 108.910 123.815 ;
        RECT 103.180 111.055 108.910 113.215 ;
        RECT 109.390 110.575 109.560 124.295 ;
        RECT 109.920 110.575 110.090 124.295 ;
        RECT 110.570 121.655 116.300 123.815 ;
        RECT 110.570 111.055 116.300 113.215 ;
        RECT 116.780 110.575 116.950 124.295 ;
        RECT 117.310 110.575 117.480 124.295 ;
        RECT 117.960 121.655 123.690 123.815 ;
        RECT 117.960 111.055 123.690 113.215 ;
        RECT 124.170 110.575 124.340 124.295 ;
        RECT 124.700 110.575 124.870 124.295 ;
        RECT 125.350 121.655 131.080 123.815 ;
        RECT 125.350 111.055 131.080 113.215 ;
        RECT 131.560 110.575 131.730 124.295 ;
        RECT 132.090 110.575 132.260 124.295 ;
        RECT 132.740 121.655 138.470 123.815 ;
        RECT 132.740 111.055 138.470 113.215 ;
        RECT 138.950 110.575 139.120 124.295 ;
        RECT 139.480 110.575 139.650 124.295 ;
        RECT 140.130 121.655 145.860 123.815 ;
        RECT 140.130 111.055 145.860 113.215 ;
        RECT 146.340 110.575 146.510 124.295 ;
        RECT 146.870 110.575 147.040 124.295 ;
        RECT 147.520 121.655 153.250 123.815 ;
        RECT 147.520 111.055 153.250 113.215 ;
        RECT 153.730 110.575 153.900 124.295 ;
        RECT 79.850 110.410 153.900 110.575 ;
        RECT 6.310 110.240 153.900 110.410 ;
        RECT 6.310 102.250 6.480 110.240 ;
        RECT 6.960 107.600 12.690 109.760 ;
        RECT 6.960 102.730 12.690 104.890 ;
        RECT 13.170 102.250 13.340 110.240 ;
        RECT 13.700 102.250 13.870 110.240 ;
        RECT 14.350 107.600 20.080 109.760 ;
        RECT 14.350 102.730 20.080 104.890 ;
        RECT 20.560 102.250 20.730 110.240 ;
        RECT 21.090 102.250 21.260 110.240 ;
        RECT 21.740 107.600 27.470 109.760 ;
        RECT 21.740 102.730 27.470 104.890 ;
        RECT 27.950 102.250 28.120 110.240 ;
        RECT 28.480 102.250 28.650 110.240 ;
        RECT 29.130 107.600 34.860 109.760 ;
        RECT 29.130 102.730 34.860 104.890 ;
        RECT 35.340 102.250 35.510 110.240 ;
        RECT 35.870 102.250 36.040 110.240 ;
        RECT 36.520 107.600 42.250 109.760 ;
        RECT 36.520 102.730 42.250 104.890 ;
        RECT 42.730 102.250 42.900 110.240 ;
        RECT 43.260 102.250 43.430 110.240 ;
        RECT 43.910 107.600 49.640 109.760 ;
        RECT 43.910 102.730 49.640 104.890 ;
        RECT 50.120 102.250 50.290 110.240 ;
        RECT 50.650 102.250 50.820 110.240 ;
        RECT 51.300 107.600 57.030 109.760 ;
        RECT 51.300 102.730 57.030 104.890 ;
        RECT 57.510 102.250 57.680 110.240 ;
        RECT 58.040 102.250 58.210 110.240 ;
        RECT 58.690 107.600 64.420 109.760 ;
        RECT 58.690 102.730 64.420 104.890 ;
        RECT 64.900 102.250 65.070 110.240 ;
        RECT 65.430 102.250 65.600 110.240 ;
        RECT 66.080 107.600 71.810 109.760 ;
        RECT 66.080 102.730 71.810 104.890 ;
        RECT 72.290 102.250 72.460 110.240 ;
        RECT 72.820 102.250 72.990 110.240 ;
        RECT 79.680 109.875 153.900 110.240 ;
        RECT 73.470 107.600 79.200 109.760 ;
        RECT 73.470 102.730 79.200 104.890 ;
        RECT 79.680 102.250 80.530 109.875 ;
        RECT 81.010 107.235 86.740 109.395 ;
        RECT 6.310 101.550 80.530 102.250 ;
        RECT 6.310 93.560 6.480 101.550 ;
        RECT 6.960 98.910 12.690 101.070 ;
        RECT 6.960 94.040 12.690 96.200 ;
        RECT 13.170 93.560 13.340 101.550 ;
        RECT 13.700 93.560 13.870 101.550 ;
        RECT 14.350 98.910 20.080 101.070 ;
        RECT 14.350 94.040 20.080 96.200 ;
        RECT 20.560 93.560 20.730 101.550 ;
        RECT 21.090 93.560 21.260 101.550 ;
        RECT 21.740 98.910 27.470 101.070 ;
        RECT 21.740 94.040 27.470 96.200 ;
        RECT 27.950 93.560 28.120 101.550 ;
        RECT 28.480 93.560 28.650 101.550 ;
        RECT 29.130 98.910 34.860 101.070 ;
        RECT 29.130 94.040 34.860 96.200 ;
        RECT 35.340 93.560 35.510 101.550 ;
        RECT 35.870 93.560 36.040 101.550 ;
        RECT 36.520 98.910 42.250 101.070 ;
        RECT 36.520 94.040 42.250 96.200 ;
        RECT 42.730 93.560 42.900 101.550 ;
        RECT 43.260 93.560 43.430 101.550 ;
        RECT 43.910 98.910 49.640 101.070 ;
        RECT 43.910 94.040 49.640 96.200 ;
        RECT 50.120 93.560 50.290 101.550 ;
        RECT 50.650 93.560 50.820 101.550 ;
        RECT 51.300 98.910 57.030 101.070 ;
        RECT 51.300 94.040 57.030 96.200 ;
        RECT 57.510 93.560 57.680 101.550 ;
        RECT 58.040 93.560 58.210 101.550 ;
        RECT 58.690 98.910 64.420 101.070 ;
        RECT 58.690 94.040 64.420 96.200 ;
        RECT 64.900 93.560 65.070 101.550 ;
        RECT 65.430 93.560 65.600 101.550 ;
        RECT 66.080 98.910 71.810 101.070 ;
        RECT 66.080 94.040 71.810 96.200 ;
        RECT 72.290 93.560 72.460 101.550 ;
        RECT 72.820 93.560 72.990 101.550 ;
        RECT 73.470 98.910 79.200 101.070 ;
        RECT 73.470 94.040 79.200 96.200 ;
        RECT 79.680 96.155 80.530 101.550 ;
        RECT 81.010 96.635 86.740 98.795 ;
        RECT 87.220 96.155 87.390 109.875 ;
        RECT 87.750 96.155 87.920 109.875 ;
        RECT 88.400 107.235 94.130 109.395 ;
        RECT 88.400 96.635 94.130 98.795 ;
        RECT 94.610 96.155 94.780 109.875 ;
        RECT 95.140 96.155 95.310 109.875 ;
        RECT 95.790 107.235 101.520 109.395 ;
        RECT 95.790 96.635 101.520 98.795 ;
        RECT 102.000 96.155 102.170 109.875 ;
        RECT 102.530 96.155 102.700 109.875 ;
        RECT 103.180 107.235 108.910 109.395 ;
        RECT 103.180 96.635 108.910 98.795 ;
        RECT 109.390 96.155 109.560 109.875 ;
        RECT 109.920 96.155 110.090 109.875 ;
        RECT 110.570 107.235 116.300 109.395 ;
        RECT 110.570 96.635 116.300 98.795 ;
        RECT 116.780 96.155 116.950 109.875 ;
        RECT 117.310 96.155 117.480 109.875 ;
        RECT 117.960 107.235 123.690 109.395 ;
        RECT 117.960 96.635 123.690 98.795 ;
        RECT 124.170 96.155 124.340 109.875 ;
        RECT 124.700 96.155 124.870 109.875 ;
        RECT 125.350 107.235 131.080 109.395 ;
        RECT 125.350 96.635 131.080 98.795 ;
        RECT 131.560 96.155 131.730 109.875 ;
        RECT 132.090 96.155 132.260 109.875 ;
        RECT 132.740 107.235 138.470 109.395 ;
        RECT 132.740 96.635 138.470 98.795 ;
        RECT 138.950 96.155 139.120 109.875 ;
        RECT 139.480 96.155 139.650 109.875 ;
        RECT 140.130 107.235 145.860 109.395 ;
        RECT 140.130 96.635 145.860 98.795 ;
        RECT 146.340 96.155 146.510 109.875 ;
        RECT 146.870 96.155 147.040 109.875 ;
        RECT 147.520 107.235 153.250 109.395 ;
        RECT 147.520 96.635 153.250 98.795 ;
        RECT 153.730 96.155 153.900 109.875 ;
        RECT 79.680 95.455 153.900 96.155 ;
        RECT 79.680 93.560 80.530 95.455 ;
        RECT 6.310 92.860 80.530 93.560 ;
        RECT 6.310 84.870 6.480 92.860 ;
        RECT 6.960 90.220 12.690 92.380 ;
        RECT 6.960 85.350 12.690 87.510 ;
        RECT 13.170 84.870 13.340 92.860 ;
        RECT 13.700 84.870 13.870 92.860 ;
        RECT 14.350 90.220 20.080 92.380 ;
        RECT 14.350 85.350 20.080 87.510 ;
        RECT 20.560 84.870 20.730 92.860 ;
        RECT 21.090 84.870 21.260 92.860 ;
        RECT 21.740 90.220 27.470 92.380 ;
        RECT 21.740 85.350 27.470 87.510 ;
        RECT 27.950 84.870 28.120 92.860 ;
        RECT 28.480 84.870 28.650 92.860 ;
        RECT 29.130 90.220 34.860 92.380 ;
        RECT 29.130 85.350 34.860 87.510 ;
        RECT 35.340 84.870 35.510 92.860 ;
        RECT 35.870 84.870 36.040 92.860 ;
        RECT 36.520 90.220 42.250 92.380 ;
        RECT 36.520 85.350 42.250 87.510 ;
        RECT 42.730 84.870 42.900 92.860 ;
        RECT 43.260 84.870 43.430 92.860 ;
        RECT 43.910 90.220 49.640 92.380 ;
        RECT 43.910 85.350 49.640 87.510 ;
        RECT 50.120 84.870 50.290 92.860 ;
        RECT 50.650 84.870 50.820 92.860 ;
        RECT 51.300 90.220 57.030 92.380 ;
        RECT 51.300 85.350 57.030 87.510 ;
        RECT 57.510 84.870 57.680 92.860 ;
        RECT 58.040 84.870 58.210 92.860 ;
        RECT 58.690 90.220 64.420 92.380 ;
        RECT 58.690 85.350 64.420 87.510 ;
        RECT 64.900 84.870 65.070 92.860 ;
        RECT 65.430 84.870 65.600 92.860 ;
        RECT 66.080 90.220 71.810 92.380 ;
        RECT 66.080 85.350 71.810 87.510 ;
        RECT 72.290 84.870 72.460 92.860 ;
        RECT 72.820 84.870 72.990 92.860 ;
        RECT 73.470 90.220 79.200 92.380 ;
        RECT 73.470 85.350 79.200 87.510 ;
        RECT 79.680 84.870 80.530 92.860 ;
        RECT 81.010 92.815 86.740 94.975 ;
        RECT 6.310 84.170 80.530 84.870 ;
        RECT 6.310 76.180 6.480 84.170 ;
        RECT 6.960 81.530 12.690 83.690 ;
        RECT 6.960 76.660 12.690 78.820 ;
        RECT 13.170 76.180 13.340 84.170 ;
        RECT 13.700 76.180 13.870 84.170 ;
        RECT 14.350 81.530 20.080 83.690 ;
        RECT 14.350 76.660 20.080 78.820 ;
        RECT 20.560 76.180 20.730 84.170 ;
        RECT 21.090 76.180 21.260 84.170 ;
        RECT 21.740 81.530 27.470 83.690 ;
        RECT 21.740 76.660 27.470 78.820 ;
        RECT 27.950 76.180 28.120 84.170 ;
        RECT 28.480 76.180 28.650 84.170 ;
        RECT 29.130 81.530 34.860 83.690 ;
        RECT 29.130 76.660 34.860 78.820 ;
        RECT 35.340 76.180 35.510 84.170 ;
        RECT 35.870 76.180 36.040 84.170 ;
        RECT 36.520 81.530 42.250 83.690 ;
        RECT 36.520 76.660 42.250 78.820 ;
        RECT 42.730 76.180 42.900 84.170 ;
        RECT 43.260 76.180 43.430 84.170 ;
        RECT 43.910 81.530 49.640 83.690 ;
        RECT 43.910 76.660 49.640 78.820 ;
        RECT 50.120 76.180 50.290 84.170 ;
        RECT 50.650 76.180 50.820 84.170 ;
        RECT 51.300 81.530 57.030 83.690 ;
        RECT 51.300 76.660 57.030 78.820 ;
        RECT 57.510 76.180 57.680 84.170 ;
        RECT 58.040 76.180 58.210 84.170 ;
        RECT 58.690 81.530 64.420 83.690 ;
        RECT 58.690 76.660 64.420 78.820 ;
        RECT 64.900 76.180 65.070 84.170 ;
        RECT 65.430 76.180 65.600 84.170 ;
        RECT 66.080 81.530 71.810 83.690 ;
        RECT 66.080 76.660 71.810 78.820 ;
        RECT 72.290 76.180 72.460 84.170 ;
        RECT 72.820 76.180 72.990 84.170 ;
        RECT 73.470 81.530 79.200 83.690 ;
        RECT 79.680 81.735 80.530 84.170 ;
        RECT 81.010 82.215 86.740 84.375 ;
        RECT 87.220 81.735 87.390 95.455 ;
        RECT 87.750 81.735 87.920 95.455 ;
        RECT 88.400 92.815 94.130 94.975 ;
        RECT 88.400 82.215 94.130 84.375 ;
        RECT 94.610 81.735 94.780 95.455 ;
        RECT 95.140 81.735 95.310 95.455 ;
        RECT 95.790 92.815 101.520 94.975 ;
        RECT 95.790 82.215 101.520 84.375 ;
        RECT 102.000 81.735 102.170 95.455 ;
        RECT 102.530 81.735 102.700 95.455 ;
        RECT 103.180 92.815 108.910 94.975 ;
        RECT 103.180 82.215 108.910 84.375 ;
        RECT 109.390 81.735 109.560 95.455 ;
        RECT 109.920 81.735 110.090 95.455 ;
        RECT 110.570 92.815 116.300 94.975 ;
        RECT 110.570 82.215 116.300 84.375 ;
        RECT 116.780 81.735 116.950 95.455 ;
        RECT 117.310 81.735 117.480 95.455 ;
        RECT 117.960 92.815 123.690 94.975 ;
        RECT 117.960 82.215 123.690 84.375 ;
        RECT 124.170 81.735 124.340 95.455 ;
        RECT 124.700 81.735 124.870 95.455 ;
        RECT 125.350 92.815 131.080 94.975 ;
        RECT 125.350 82.215 131.080 84.375 ;
        RECT 131.560 81.735 131.730 95.455 ;
        RECT 132.090 81.735 132.260 95.455 ;
        RECT 132.740 92.815 138.470 94.975 ;
        RECT 132.740 82.215 138.470 84.375 ;
        RECT 138.950 81.735 139.120 95.455 ;
        RECT 139.480 81.735 139.650 95.455 ;
        RECT 140.130 92.815 145.860 94.975 ;
        RECT 140.130 82.215 145.860 84.375 ;
        RECT 146.340 81.735 146.510 95.455 ;
        RECT 146.870 81.735 147.040 95.455 ;
        RECT 147.520 92.815 153.250 94.975 ;
        RECT 147.520 82.215 153.250 84.375 ;
        RECT 153.730 81.735 153.900 95.455 ;
        RECT 79.680 81.035 153.900 81.735 ;
        RECT 73.470 76.660 79.200 78.820 ;
        RECT 79.680 76.180 80.530 81.035 ;
        RECT 81.010 78.395 86.740 80.555 ;
        RECT 6.310 75.480 80.530 76.180 ;
        RECT 6.310 67.490 6.480 75.480 ;
        RECT 6.960 72.840 12.690 75.000 ;
        RECT 6.960 67.970 12.690 70.130 ;
        RECT 13.170 67.490 13.340 75.480 ;
        RECT 13.700 67.490 13.870 75.480 ;
        RECT 14.350 72.840 20.080 75.000 ;
        RECT 14.350 67.970 20.080 70.130 ;
        RECT 20.560 67.490 20.730 75.480 ;
        RECT 21.090 67.490 21.260 75.480 ;
        RECT 21.740 72.840 27.470 75.000 ;
        RECT 21.740 67.970 27.470 70.130 ;
        RECT 27.950 67.490 28.120 75.480 ;
        RECT 28.480 67.490 28.650 75.480 ;
        RECT 29.130 72.840 34.860 75.000 ;
        RECT 29.130 67.970 34.860 70.130 ;
        RECT 35.340 67.490 35.510 75.480 ;
        RECT 35.870 67.490 36.040 75.480 ;
        RECT 36.520 72.840 42.250 75.000 ;
        RECT 36.520 67.970 42.250 70.130 ;
        RECT 42.730 67.490 42.900 75.480 ;
        RECT 43.260 67.490 43.430 75.480 ;
        RECT 43.910 72.840 49.640 75.000 ;
        RECT 43.910 67.970 49.640 70.130 ;
        RECT 50.120 67.490 50.290 75.480 ;
        RECT 50.650 67.490 50.820 75.480 ;
        RECT 51.300 72.840 57.030 75.000 ;
        RECT 51.300 67.970 57.030 70.130 ;
        RECT 57.510 67.490 57.680 75.480 ;
        RECT 58.040 67.490 58.210 75.480 ;
        RECT 58.690 72.840 64.420 75.000 ;
        RECT 58.690 67.970 64.420 70.130 ;
        RECT 64.900 67.490 65.070 75.480 ;
        RECT 65.430 67.490 65.600 75.480 ;
        RECT 66.080 72.840 71.810 75.000 ;
        RECT 66.080 67.970 71.810 70.130 ;
        RECT 72.290 67.490 72.460 75.480 ;
        RECT 72.820 67.490 72.990 75.480 ;
        RECT 73.470 72.840 79.200 75.000 ;
        RECT 73.470 67.970 79.200 70.130 ;
        RECT 79.680 67.490 80.530 75.480 ;
        RECT 81.010 67.795 86.740 69.955 ;
        RECT 6.310 67.315 80.530 67.490 ;
        RECT 87.220 67.315 87.390 81.035 ;
        RECT 87.750 67.315 87.920 81.035 ;
        RECT 88.400 78.395 94.130 80.555 ;
        RECT 88.400 67.795 94.130 69.955 ;
        RECT 94.610 67.315 94.780 81.035 ;
        RECT 95.140 67.315 95.310 81.035 ;
        RECT 95.790 78.395 101.520 80.555 ;
        RECT 95.790 67.795 101.520 69.955 ;
        RECT 102.000 67.315 102.170 81.035 ;
        RECT 102.530 67.315 102.700 81.035 ;
        RECT 103.180 78.395 108.910 80.555 ;
        RECT 103.180 67.795 108.910 69.955 ;
        RECT 109.390 67.315 109.560 81.035 ;
        RECT 109.920 67.315 110.090 81.035 ;
        RECT 110.570 78.395 116.300 80.555 ;
        RECT 110.570 67.795 116.300 69.955 ;
        RECT 116.780 67.315 116.950 81.035 ;
        RECT 117.310 67.315 117.480 81.035 ;
        RECT 117.960 78.395 123.690 80.555 ;
        RECT 117.960 67.795 123.690 69.955 ;
        RECT 124.170 67.315 124.340 81.035 ;
        RECT 124.700 67.315 124.870 81.035 ;
        RECT 125.350 78.395 131.080 80.555 ;
        RECT 125.350 67.795 131.080 69.955 ;
        RECT 131.560 67.315 131.730 81.035 ;
        RECT 132.090 67.315 132.260 81.035 ;
        RECT 132.740 78.395 138.470 80.555 ;
        RECT 132.740 67.795 138.470 69.955 ;
        RECT 138.950 67.315 139.120 81.035 ;
        RECT 139.480 67.315 139.650 81.035 ;
        RECT 140.130 78.395 145.860 80.555 ;
        RECT 140.130 67.795 145.860 69.955 ;
        RECT 146.340 67.315 146.510 81.035 ;
        RECT 146.870 67.315 147.040 81.035 ;
        RECT 147.520 78.395 153.250 80.555 ;
        RECT 147.520 67.795 153.250 69.955 ;
        RECT 153.730 67.315 153.900 81.035 ;
        RECT 6.310 66.790 153.900 67.315 ;
        RECT 6.310 58.800 6.480 66.790 ;
        RECT 6.960 64.150 12.690 66.310 ;
        RECT 6.960 59.280 12.690 61.440 ;
        RECT 13.170 58.800 13.340 66.790 ;
        RECT 13.700 58.800 13.870 66.790 ;
        RECT 14.350 64.150 20.080 66.310 ;
        RECT 14.350 59.280 20.080 61.440 ;
        RECT 20.560 58.800 20.730 66.790 ;
        RECT 21.090 58.800 21.260 66.790 ;
        RECT 21.740 64.150 27.470 66.310 ;
        RECT 21.740 59.280 27.470 61.440 ;
        RECT 27.950 58.800 28.120 66.790 ;
        RECT 28.480 58.800 28.650 66.790 ;
        RECT 29.130 64.150 34.860 66.310 ;
        RECT 29.130 59.280 34.860 61.440 ;
        RECT 35.340 58.800 35.510 66.790 ;
        RECT 35.870 58.800 36.040 66.790 ;
        RECT 36.520 64.150 42.250 66.310 ;
        RECT 36.520 59.280 42.250 61.440 ;
        RECT 42.730 58.800 42.900 66.790 ;
        RECT 43.260 58.800 43.430 66.790 ;
        RECT 43.910 64.150 49.640 66.310 ;
        RECT 43.910 59.280 49.640 61.440 ;
        RECT 50.120 58.800 50.290 66.790 ;
        RECT 50.650 58.800 50.820 66.790 ;
        RECT 51.300 64.150 57.030 66.310 ;
        RECT 51.300 59.280 57.030 61.440 ;
        RECT 57.510 58.800 57.680 66.790 ;
        RECT 58.040 58.800 58.210 66.790 ;
        RECT 58.690 64.150 64.420 66.310 ;
        RECT 58.690 59.280 64.420 61.440 ;
        RECT 64.900 58.800 65.070 66.790 ;
        RECT 65.430 58.800 65.600 66.790 ;
        RECT 66.080 64.150 71.810 66.310 ;
        RECT 66.080 59.280 71.810 61.440 ;
        RECT 72.290 58.800 72.460 66.790 ;
        RECT 72.820 58.800 72.990 66.790 ;
        RECT 79.680 66.615 153.900 66.790 ;
        RECT 73.470 64.150 79.200 66.310 ;
        RECT 73.470 59.280 79.200 61.440 ;
        RECT 79.680 58.800 80.530 66.615 ;
        RECT 81.010 63.975 86.740 66.135 ;
        RECT 6.310 58.100 80.530 58.800 ;
        RECT 6.310 50.110 6.480 58.100 ;
        RECT 6.960 55.460 12.690 57.620 ;
        RECT 6.960 50.590 12.690 52.750 ;
        RECT 13.170 50.110 13.340 58.100 ;
        RECT 13.700 50.110 13.870 58.100 ;
        RECT 14.350 55.460 20.080 57.620 ;
        RECT 14.350 50.590 20.080 52.750 ;
        RECT 20.560 50.110 20.730 58.100 ;
        RECT 21.090 50.110 21.260 58.100 ;
        RECT 21.740 55.460 27.470 57.620 ;
        RECT 21.740 50.590 27.470 52.750 ;
        RECT 27.950 50.110 28.120 58.100 ;
        RECT 28.480 50.110 28.650 58.100 ;
        RECT 29.130 55.460 34.860 57.620 ;
        RECT 29.130 50.590 34.860 52.750 ;
        RECT 35.340 50.110 35.510 58.100 ;
        RECT 35.870 50.110 36.040 58.100 ;
        RECT 36.520 55.460 42.250 57.620 ;
        RECT 36.520 50.590 42.250 52.750 ;
        RECT 42.730 50.110 42.900 58.100 ;
        RECT 43.260 50.110 43.430 58.100 ;
        RECT 43.910 55.460 49.640 57.620 ;
        RECT 43.910 50.590 49.640 52.750 ;
        RECT 50.120 50.110 50.290 58.100 ;
        RECT 50.650 50.110 50.820 58.100 ;
        RECT 51.300 55.460 57.030 57.620 ;
        RECT 51.300 50.590 57.030 52.750 ;
        RECT 57.510 50.110 57.680 58.100 ;
        RECT 58.040 50.110 58.210 58.100 ;
        RECT 58.690 55.460 64.420 57.620 ;
        RECT 58.690 50.590 64.420 52.750 ;
        RECT 64.900 50.110 65.070 58.100 ;
        RECT 65.430 50.110 65.600 58.100 ;
        RECT 66.080 55.460 71.810 57.620 ;
        RECT 66.080 50.590 71.810 52.750 ;
        RECT 72.290 50.110 72.460 58.100 ;
        RECT 72.820 50.110 72.990 58.100 ;
        RECT 73.470 55.460 79.200 57.620 ;
        RECT 79.680 52.895 80.530 58.100 ;
        RECT 81.010 53.375 86.740 55.535 ;
        RECT 87.220 52.895 87.390 66.615 ;
        RECT 87.750 52.895 87.920 66.615 ;
        RECT 88.400 63.975 94.130 66.135 ;
        RECT 88.400 53.375 94.130 55.535 ;
        RECT 94.610 52.895 94.780 66.615 ;
        RECT 95.140 52.895 95.310 66.615 ;
        RECT 95.790 63.975 101.520 66.135 ;
        RECT 95.790 53.375 101.520 55.535 ;
        RECT 102.000 52.895 102.170 66.615 ;
        RECT 102.530 52.895 102.700 66.615 ;
        RECT 103.180 63.975 108.910 66.135 ;
        RECT 103.180 53.375 108.910 55.535 ;
        RECT 109.390 52.895 109.560 66.615 ;
        RECT 109.920 52.895 110.090 66.615 ;
        RECT 110.570 63.975 116.300 66.135 ;
        RECT 110.570 53.375 116.300 55.535 ;
        RECT 116.780 52.895 116.950 66.615 ;
        RECT 117.310 52.895 117.480 66.615 ;
        RECT 117.960 63.975 123.690 66.135 ;
        RECT 117.960 53.375 123.690 55.535 ;
        RECT 124.170 52.895 124.340 66.615 ;
        RECT 124.700 52.895 124.870 66.615 ;
        RECT 125.350 63.975 131.080 66.135 ;
        RECT 125.350 53.375 131.080 55.535 ;
        RECT 131.560 52.895 131.730 66.615 ;
        RECT 132.090 52.895 132.260 66.615 ;
        RECT 132.740 63.975 138.470 66.135 ;
        RECT 132.740 53.375 138.470 55.535 ;
        RECT 138.950 52.895 139.120 66.615 ;
        RECT 139.480 52.895 139.650 66.615 ;
        RECT 140.130 63.975 145.860 66.135 ;
        RECT 140.130 53.375 145.860 55.535 ;
        RECT 146.340 52.895 146.510 66.615 ;
        RECT 146.870 52.895 147.040 66.615 ;
        RECT 147.520 63.975 153.250 66.135 ;
        RECT 147.520 53.375 153.250 55.535 ;
        RECT 153.730 52.895 153.900 66.615 ;
        RECT 73.470 50.590 79.200 52.750 ;
        RECT 79.680 52.195 153.900 52.895 ;
        RECT 79.680 50.110 80.530 52.195 ;
        RECT 6.310 49.410 80.530 50.110 ;
        RECT 81.010 49.555 86.740 51.715 ;
        RECT 6.310 41.420 6.480 49.410 ;
        RECT 6.960 46.770 12.690 48.930 ;
        RECT 6.960 41.900 12.690 44.060 ;
        RECT 13.170 41.420 13.340 49.410 ;
        RECT 13.700 41.420 13.870 49.410 ;
        RECT 14.350 46.770 20.080 48.930 ;
        RECT 14.350 41.900 20.080 44.060 ;
        RECT 20.560 41.420 20.730 49.410 ;
        RECT 21.090 41.420 21.260 49.410 ;
        RECT 21.740 46.770 27.470 48.930 ;
        RECT 21.740 41.900 27.470 44.060 ;
        RECT 27.950 41.420 28.120 49.410 ;
        RECT 28.480 41.420 28.650 49.410 ;
        RECT 29.130 46.770 34.860 48.930 ;
        RECT 29.130 41.900 34.860 44.060 ;
        RECT 35.340 41.420 35.510 49.410 ;
        RECT 35.870 41.420 36.040 49.410 ;
        RECT 36.520 46.770 42.250 48.930 ;
        RECT 36.520 41.900 42.250 44.060 ;
        RECT 42.730 41.420 42.900 49.410 ;
        RECT 43.260 41.420 43.430 49.410 ;
        RECT 43.910 46.770 49.640 48.930 ;
        RECT 43.910 41.900 49.640 44.060 ;
        RECT 50.120 41.420 50.290 49.410 ;
        RECT 50.650 41.420 50.820 49.410 ;
        RECT 51.300 46.770 57.030 48.930 ;
        RECT 51.300 41.900 57.030 44.060 ;
        RECT 57.510 41.420 57.680 49.410 ;
        RECT 58.040 41.420 58.210 49.410 ;
        RECT 58.690 46.770 64.420 48.930 ;
        RECT 58.690 41.900 64.420 44.060 ;
        RECT 64.900 41.420 65.070 49.410 ;
        RECT 65.430 41.420 65.600 49.410 ;
        RECT 66.080 46.770 71.810 48.930 ;
        RECT 66.080 41.900 71.810 44.060 ;
        RECT 72.290 41.420 72.460 49.410 ;
        RECT 72.820 41.420 72.990 49.410 ;
        RECT 73.470 46.770 79.200 48.930 ;
        RECT 73.470 41.900 79.200 44.060 ;
        RECT 79.680 41.420 80.530 49.410 ;
        RECT 6.310 40.720 80.530 41.420 ;
        RECT 6.310 32.730 6.480 40.720 ;
        RECT 6.960 38.080 12.690 40.240 ;
        RECT 6.960 33.210 12.690 35.370 ;
        RECT 13.170 32.730 13.340 40.720 ;
        RECT 13.700 32.730 13.870 40.720 ;
        RECT 14.350 38.080 20.080 40.240 ;
        RECT 14.350 33.210 20.080 35.370 ;
        RECT 20.560 32.730 20.730 40.720 ;
        RECT 21.090 32.730 21.260 40.720 ;
        RECT 21.740 38.080 27.470 40.240 ;
        RECT 21.740 33.210 27.470 35.370 ;
        RECT 27.950 32.730 28.120 40.720 ;
        RECT 28.480 32.730 28.650 40.720 ;
        RECT 29.130 38.080 34.860 40.240 ;
        RECT 29.130 33.210 34.860 35.370 ;
        RECT 35.340 32.730 35.510 40.720 ;
        RECT 35.870 32.730 36.040 40.720 ;
        RECT 36.520 38.080 42.250 40.240 ;
        RECT 36.520 33.210 42.250 35.370 ;
        RECT 42.730 32.730 42.900 40.720 ;
        RECT 43.260 32.730 43.430 40.720 ;
        RECT 43.910 38.080 49.640 40.240 ;
        RECT 43.910 33.210 49.640 35.370 ;
        RECT 50.120 32.730 50.290 40.720 ;
        RECT 50.650 32.730 50.820 40.720 ;
        RECT 51.300 38.080 57.030 40.240 ;
        RECT 51.300 33.210 57.030 35.370 ;
        RECT 57.510 32.730 57.680 40.720 ;
        RECT 58.040 32.730 58.210 40.720 ;
        RECT 58.690 38.080 64.420 40.240 ;
        RECT 58.690 33.210 64.420 35.370 ;
        RECT 64.900 32.730 65.070 40.720 ;
        RECT 65.430 32.730 65.600 40.720 ;
        RECT 66.080 38.080 71.810 40.240 ;
        RECT 66.080 33.210 71.810 35.370 ;
        RECT 72.290 32.730 72.460 40.720 ;
        RECT 72.820 32.730 72.990 40.720 ;
        RECT 73.470 38.080 79.200 40.240 ;
        RECT 79.680 38.475 80.530 40.720 ;
        RECT 81.010 38.955 86.740 41.115 ;
        RECT 87.220 38.475 87.390 52.195 ;
        RECT 87.750 38.475 87.920 52.195 ;
        RECT 88.400 49.555 94.130 51.715 ;
        RECT 88.400 38.955 94.130 41.115 ;
        RECT 94.610 38.475 94.780 52.195 ;
        RECT 95.140 38.475 95.310 52.195 ;
        RECT 95.790 49.555 101.520 51.715 ;
        RECT 95.790 38.955 101.520 41.115 ;
        RECT 102.000 38.475 102.170 52.195 ;
        RECT 102.530 38.475 102.700 52.195 ;
        RECT 103.180 49.555 108.910 51.715 ;
        RECT 103.180 38.955 108.910 41.115 ;
        RECT 109.390 38.475 109.560 52.195 ;
        RECT 109.920 38.475 110.090 52.195 ;
        RECT 110.570 49.555 116.300 51.715 ;
        RECT 110.570 38.955 116.300 41.115 ;
        RECT 116.780 38.475 116.950 52.195 ;
        RECT 117.310 38.475 117.480 52.195 ;
        RECT 117.960 49.555 123.690 51.715 ;
        RECT 117.960 38.955 123.690 41.115 ;
        RECT 124.170 38.475 124.340 52.195 ;
        RECT 124.700 38.475 124.870 52.195 ;
        RECT 125.350 49.555 131.080 51.715 ;
        RECT 125.350 38.955 131.080 41.115 ;
        RECT 131.560 38.475 131.730 52.195 ;
        RECT 132.090 38.475 132.260 52.195 ;
        RECT 132.740 49.555 138.470 51.715 ;
        RECT 132.740 38.955 138.470 41.115 ;
        RECT 138.950 38.475 139.120 52.195 ;
        RECT 139.480 38.475 139.650 52.195 ;
        RECT 140.130 49.555 145.860 51.715 ;
        RECT 140.130 38.955 145.860 41.115 ;
        RECT 146.340 38.475 146.510 52.195 ;
        RECT 146.870 38.475 147.040 52.195 ;
        RECT 147.520 49.555 153.250 51.715 ;
        RECT 147.520 38.955 153.250 41.115 ;
        RECT 153.730 38.475 153.900 52.195 ;
        RECT 79.680 37.775 153.900 38.475 ;
        RECT 73.470 33.210 79.200 35.370 ;
        RECT 79.680 32.730 80.530 37.775 ;
        RECT 81.010 35.135 86.740 37.295 ;
        RECT 6.310 32.030 80.530 32.730 ;
        RECT 6.310 24.040 6.480 32.030 ;
        RECT 6.960 29.390 12.690 31.550 ;
        RECT 6.960 24.520 12.690 26.680 ;
        RECT 13.170 24.040 13.340 32.030 ;
        RECT 13.700 24.040 13.870 32.030 ;
        RECT 14.350 29.390 20.080 31.550 ;
        RECT 14.350 24.520 20.080 26.680 ;
        RECT 20.560 24.040 20.730 32.030 ;
        RECT 21.090 24.040 21.260 32.030 ;
        RECT 21.740 29.390 27.470 31.550 ;
        RECT 21.740 24.520 27.470 26.680 ;
        RECT 27.950 24.040 28.120 32.030 ;
        RECT 28.480 24.040 28.650 32.030 ;
        RECT 29.130 29.390 34.860 31.550 ;
        RECT 29.130 24.520 34.860 26.680 ;
        RECT 35.340 24.040 35.510 32.030 ;
        RECT 35.870 24.040 36.040 32.030 ;
        RECT 36.520 29.390 42.250 31.550 ;
        RECT 36.520 24.520 42.250 26.680 ;
        RECT 42.730 24.040 42.900 32.030 ;
        RECT 43.260 24.040 43.430 32.030 ;
        RECT 43.910 29.390 49.640 31.550 ;
        RECT 43.910 24.520 49.640 26.680 ;
        RECT 50.120 24.040 50.290 32.030 ;
        RECT 50.650 24.040 50.820 32.030 ;
        RECT 51.300 29.390 57.030 31.550 ;
        RECT 51.300 24.520 57.030 26.680 ;
        RECT 57.510 24.040 57.680 32.030 ;
        RECT 58.040 24.040 58.210 32.030 ;
        RECT 58.690 29.390 64.420 31.550 ;
        RECT 58.690 24.520 64.420 26.680 ;
        RECT 64.900 24.040 65.070 32.030 ;
        RECT 65.430 24.040 65.600 32.030 ;
        RECT 66.080 29.390 71.810 31.550 ;
        RECT 66.080 24.520 71.810 26.680 ;
        RECT 72.290 24.040 72.460 32.030 ;
        RECT 72.820 24.040 72.990 32.030 ;
        RECT 73.470 29.390 79.200 31.550 ;
        RECT 73.470 24.520 79.200 26.680 ;
        RECT 79.680 24.055 80.530 32.030 ;
        RECT 81.010 24.535 86.740 26.695 ;
        RECT 87.220 24.055 87.390 37.775 ;
        RECT 87.750 24.055 87.920 37.775 ;
        RECT 88.400 35.135 94.130 37.295 ;
        RECT 88.400 24.535 94.130 26.695 ;
        RECT 94.610 24.055 94.780 37.775 ;
        RECT 95.140 24.055 95.310 37.775 ;
        RECT 95.790 35.135 101.520 37.295 ;
        RECT 95.790 24.535 101.520 26.695 ;
        RECT 102.000 24.055 102.170 37.775 ;
        RECT 102.530 24.055 102.700 37.775 ;
        RECT 103.180 35.135 108.910 37.295 ;
        RECT 103.180 24.535 108.910 26.695 ;
        RECT 109.390 24.055 109.560 37.775 ;
        RECT 109.920 24.055 110.090 37.775 ;
        RECT 110.570 35.135 116.300 37.295 ;
        RECT 110.570 24.535 116.300 26.695 ;
        RECT 116.780 24.055 116.950 37.775 ;
        RECT 117.310 24.055 117.480 37.775 ;
        RECT 117.960 35.135 123.690 37.295 ;
        RECT 117.960 24.535 123.690 26.695 ;
        RECT 124.170 24.055 124.340 37.775 ;
        RECT 124.700 24.055 124.870 37.775 ;
        RECT 125.350 35.135 131.080 37.295 ;
        RECT 125.350 24.535 131.080 26.695 ;
        RECT 131.560 24.055 131.730 37.775 ;
        RECT 132.090 24.055 132.260 37.775 ;
        RECT 132.740 35.135 138.470 37.295 ;
        RECT 132.740 24.535 138.470 26.695 ;
        RECT 138.950 24.055 139.120 37.775 ;
        RECT 139.480 24.055 139.650 37.775 ;
        RECT 140.130 35.135 145.860 37.295 ;
        RECT 140.130 24.535 145.860 26.695 ;
        RECT 146.340 24.055 146.510 37.775 ;
        RECT 146.870 24.055 147.040 37.775 ;
        RECT 147.520 35.135 153.250 37.295 ;
        RECT 147.520 24.535 153.250 26.695 ;
        RECT 153.730 24.055 153.900 37.775 ;
        RECT 79.680 24.040 153.900 24.055 ;
        RECT 6.310 21.435 153.900 24.040 ;
        RECT 6.310 19.050 102.795 21.435 ;
        RECT 114.635 21.320 153.900 21.435 ;
        RECT 6.310 5.330 11.110 19.050 ;
        RECT 11.590 16.410 17.320 18.570 ;
        RECT 11.590 5.810 17.320 7.970 ;
        RECT 17.800 5.330 17.970 19.050 ;
        RECT 6.310 5.270 17.970 5.330 ;
        RECT 18.330 5.330 18.500 19.050 ;
        RECT 18.980 16.410 24.710 18.570 ;
        RECT 18.980 5.810 24.710 7.970 ;
        RECT 25.190 5.330 25.360 19.050 ;
        RECT 18.330 5.270 25.360 5.330 ;
        RECT 25.720 5.330 25.890 19.050 ;
        RECT 26.370 16.410 32.100 18.570 ;
        RECT 26.370 5.810 32.100 7.970 ;
        RECT 32.580 5.330 32.750 19.050 ;
        RECT 25.720 5.270 32.750 5.330 ;
        RECT 33.110 5.330 33.280 19.050 ;
        RECT 33.760 16.410 39.490 18.570 ;
        RECT 33.760 5.810 39.490 7.970 ;
        RECT 39.970 5.330 40.140 19.050 ;
        RECT 33.110 5.270 40.140 5.330 ;
        RECT 40.500 5.330 40.670 19.050 ;
        RECT 41.150 16.410 46.880 18.570 ;
        RECT 41.150 5.810 46.880 7.970 ;
        RECT 47.360 5.330 47.530 19.050 ;
        RECT 40.500 5.270 47.530 5.330 ;
        RECT 47.890 5.330 48.060 19.050 ;
        RECT 48.540 16.410 54.270 18.570 ;
        RECT 48.540 5.810 54.270 7.970 ;
        RECT 54.750 5.330 54.920 19.050 ;
        RECT 47.890 5.270 54.920 5.330 ;
        RECT 55.280 5.330 55.450 19.050 ;
        RECT 55.930 16.410 61.660 18.570 ;
        RECT 55.930 5.810 61.660 7.970 ;
        RECT 62.140 5.330 62.310 19.050 ;
        RECT 55.280 5.270 62.310 5.330 ;
        RECT 62.670 5.330 62.840 19.050 ;
        RECT 63.320 16.410 69.050 18.570 ;
        RECT 63.320 5.810 69.050 7.970 ;
        RECT 69.530 5.330 69.700 19.050 ;
        RECT 62.670 5.270 69.700 5.330 ;
        RECT 70.060 5.330 70.230 19.050 ;
        RECT 70.710 16.410 76.440 18.570 ;
        RECT 70.710 5.810 76.440 7.970 ;
        RECT 76.920 5.330 77.090 19.050 ;
        RECT 70.060 5.270 77.090 5.330 ;
        RECT 77.450 5.330 77.620 19.050 ;
        RECT 78.100 16.410 83.830 18.570 ;
        RECT 84.310 18.325 102.795 19.050 ;
        RECT 78.100 5.810 83.830 7.970 ;
        RECT 84.310 5.330 90.955 18.325 ;
        RECT 91.435 15.685 97.165 17.845 ;
        RECT 97.645 12.475 102.795 18.325 ;
        RECT 103.225 19.100 105.325 19.680 ;
        RECT 103.225 16.610 103.395 19.100 ;
        RECT 104.025 18.590 104.525 18.760 ;
        RECT 103.795 17.335 103.965 18.375 ;
        RECT 104.585 17.335 104.755 18.375 ;
        RECT 104.025 16.950 104.525 17.120 ;
        RECT 105.155 16.610 105.325 19.100 ;
        RECT 103.225 16.440 105.325 16.610 ;
        RECT 106.185 19.100 114.205 19.680 ;
        RECT 106.185 16.610 106.355 19.100 ;
        RECT 106.985 18.590 107.485 18.760 ;
        RECT 106.755 17.335 106.925 18.375 ;
        RECT 107.545 17.335 107.715 18.375 ;
        RECT 106.985 16.950 107.485 17.120 ;
        RECT 108.115 16.610 108.285 19.100 ;
        RECT 106.185 16.440 108.285 16.610 ;
        RECT 109.145 16.610 109.315 19.100 ;
        RECT 109.945 18.590 110.445 18.760 ;
        RECT 109.715 17.335 109.885 18.375 ;
        RECT 110.505 17.335 110.675 18.375 ;
        RECT 109.945 16.950 110.445 17.120 ;
        RECT 111.075 16.610 111.245 19.100 ;
        RECT 109.145 16.440 111.245 16.610 ;
        RECT 112.105 16.610 112.275 19.100 ;
        RECT 112.905 18.590 113.405 18.760 ;
        RECT 112.675 17.335 112.845 18.375 ;
        RECT 113.465 17.335 113.635 18.375 ;
        RECT 112.905 16.950 113.405 17.120 ;
        RECT 114.035 16.610 114.205 19.100 ;
        RECT 112.105 16.440 114.205 16.610 ;
        RECT 114.635 16.975 144.420 21.320 ;
        RECT 102.975 15.225 105.575 15.395 ;
        RECT 102.975 12.825 103.145 15.225 ;
        RECT 103.775 14.715 104.775 14.885 ;
        RECT 103.545 13.505 103.715 14.545 ;
        RECT 104.835 13.505 105.005 14.545 ;
        RECT 103.775 13.165 104.775 13.335 ;
        RECT 105.405 12.825 105.575 15.225 ;
        RECT 102.975 12.475 105.575 12.825 ;
        RECT 105.935 15.225 108.535 15.395 ;
        RECT 105.935 12.825 106.105 15.225 ;
        RECT 106.735 14.715 107.735 14.885 ;
        RECT 106.505 13.505 106.675 14.545 ;
        RECT 107.795 13.505 107.965 14.545 ;
        RECT 106.735 13.165 107.735 13.335 ;
        RECT 108.365 12.825 108.535 15.225 ;
        RECT 108.895 15.225 111.495 15.395 ;
        RECT 108.895 12.825 109.065 15.225 ;
        RECT 109.695 14.715 110.695 14.885 ;
        RECT 109.465 13.505 109.635 14.545 ;
        RECT 110.755 13.505 110.925 14.545 ;
        RECT 109.695 13.165 110.695 13.335 ;
        RECT 111.325 12.825 111.495 15.225 ;
        RECT 111.855 15.225 114.455 15.395 ;
        RECT 111.855 12.825 112.025 15.225 ;
        RECT 112.655 14.715 113.655 14.885 ;
        RECT 112.425 13.505 112.595 14.545 ;
        RECT 113.715 13.505 113.885 14.545 ;
        RECT 112.655 13.165 113.655 13.335 ;
        RECT 114.285 12.825 114.455 15.225 ;
        RECT 105.935 12.475 114.455 12.825 ;
        RECT 114.635 12.475 129.595 16.975 ;
        RECT 130.075 14.335 135.805 16.495 ;
        RECT 97.645 11.785 129.595 12.475 ;
        RECT 77.450 5.270 90.955 5.330 ;
        RECT 6.310 4.605 90.955 5.270 ;
        RECT 91.435 5.085 97.165 7.245 ;
        RECT 97.645 4.605 102.795 11.785 ;
        RECT 102.975 11.435 105.575 11.785 ;
        RECT 102.975 9.035 103.145 11.435 ;
        RECT 103.775 10.925 104.775 11.095 ;
        RECT 103.545 9.715 103.715 10.755 ;
        RECT 104.835 9.715 105.005 10.755 ;
        RECT 103.775 9.375 104.775 9.545 ;
        RECT 105.405 9.035 105.575 11.435 ;
        RECT 102.975 8.865 105.575 9.035 ;
        RECT 105.935 11.435 114.455 11.785 ;
        RECT 105.935 9.035 106.105 11.435 ;
        RECT 106.735 10.925 107.735 11.095 ;
        RECT 106.505 9.715 106.675 10.755 ;
        RECT 107.795 9.715 107.965 10.755 ;
        RECT 106.735 9.375 107.735 9.545 ;
        RECT 108.365 9.035 108.535 11.435 ;
        RECT 105.935 8.865 108.535 9.035 ;
        RECT 108.895 9.035 109.065 11.435 ;
        RECT 109.695 10.925 110.695 11.095 ;
        RECT 109.465 9.715 109.635 10.755 ;
        RECT 110.755 9.715 110.925 10.755 ;
        RECT 109.695 9.375 110.695 9.545 ;
        RECT 111.325 9.035 111.495 11.435 ;
        RECT 108.895 8.865 111.495 9.035 ;
        RECT 111.855 9.035 112.025 11.435 ;
        RECT 112.655 10.925 113.655 11.095 ;
        RECT 112.425 9.715 112.595 10.755 ;
        RECT 113.715 9.715 113.885 10.755 ;
        RECT 112.655 9.375 113.655 9.545 ;
        RECT 114.285 9.035 114.455 11.435 ;
        RECT 111.855 8.865 114.455 9.035 ;
        RECT 6.310 3.910 102.795 4.605 ;
        RECT 103.225 7.650 105.325 7.820 ;
        RECT 103.225 5.160 103.395 7.650 ;
        RECT 104.025 7.140 104.525 7.310 ;
        RECT 103.795 5.885 103.965 6.925 ;
        RECT 104.585 5.885 104.755 6.925 ;
        RECT 104.025 5.500 104.525 5.670 ;
        RECT 105.155 5.160 105.325 7.650 ;
        RECT 103.225 4.580 105.325 5.160 ;
        RECT 106.185 7.650 108.285 7.820 ;
        RECT 106.185 5.160 106.355 7.650 ;
        RECT 106.985 7.140 107.485 7.310 ;
        RECT 106.755 5.885 106.925 6.925 ;
        RECT 107.545 5.885 107.715 6.925 ;
        RECT 106.985 5.500 107.485 5.670 ;
        RECT 108.115 5.160 108.285 7.650 ;
        RECT 109.145 7.650 111.245 7.820 ;
        RECT 109.145 5.160 109.315 7.650 ;
        RECT 109.945 7.140 110.445 7.310 ;
        RECT 109.715 5.885 109.885 6.925 ;
        RECT 110.505 5.885 110.675 6.925 ;
        RECT 109.945 5.500 110.445 5.670 ;
        RECT 111.075 5.160 111.245 7.650 ;
        RECT 112.105 7.650 114.205 7.820 ;
        RECT 112.105 5.160 112.275 7.650 ;
        RECT 112.905 7.140 113.405 7.310 ;
        RECT 112.675 5.885 112.845 6.925 ;
        RECT 113.465 5.885 113.635 6.925 ;
        RECT 112.905 5.500 113.405 5.670 ;
        RECT 114.035 5.160 114.205 7.650 ;
        RECT 106.185 4.580 114.205 5.160 ;
        RECT 114.635 3.910 129.595 11.785 ;
        RECT 136.285 7.650 144.420 16.975 ;
        RECT 144.600 19.970 149.860 20.550 ;
        RECT 144.600 14.480 144.770 19.970 ;
        RECT 145.170 15.205 145.340 19.245 ;
        RECT 145.960 15.205 146.130 19.245 ;
        RECT 146.750 15.205 146.920 19.245 ;
        RECT 147.540 15.205 147.710 19.245 ;
        RECT 148.330 15.205 148.500 19.245 ;
        RECT 149.120 15.205 149.290 19.245 ;
        RECT 145.400 14.820 145.900 14.990 ;
        RECT 146.190 14.820 146.690 14.990 ;
        RECT 146.980 14.820 147.480 14.990 ;
        RECT 147.770 14.820 148.270 14.990 ;
        RECT 148.560 14.820 149.060 14.990 ;
        RECT 149.690 14.480 149.860 19.970 ;
        RECT 144.600 14.310 149.860 14.480 ;
        RECT 144.600 13.095 149.860 13.265 ;
        RECT 144.600 7.695 144.770 13.095 ;
        RECT 145.400 12.585 145.900 12.755 ;
        RECT 146.190 12.585 146.690 12.755 ;
        RECT 146.980 12.585 147.480 12.755 ;
        RECT 147.770 12.585 148.270 12.755 ;
        RECT 148.560 12.585 149.060 12.755 ;
        RECT 145.170 8.375 145.340 12.415 ;
        RECT 145.960 8.375 146.130 12.415 ;
        RECT 146.750 8.375 146.920 12.415 ;
        RECT 147.540 8.375 147.710 12.415 ;
        RECT 148.330 8.375 148.500 12.415 ;
        RECT 149.120 8.375 149.290 12.415 ;
        RECT 149.690 7.695 149.860 13.095 ;
        RECT 144.600 7.650 149.860 7.695 ;
        RECT 150.040 7.650 153.900 21.320 ;
        RECT 6.310 3.255 129.595 3.910 ;
        RECT 130.075 3.735 135.805 5.895 ;
        RECT 136.285 3.255 153.900 7.650 ;
        RECT 6.310 2.025 153.900 3.255 ;
      LAYER met1 ;
        RECT 81.010 164.915 94.130 167.075 ;
        RECT 95.790 164.915 108.910 167.075 ;
        RECT 110.570 164.915 123.690 167.075 ;
        RECT 125.350 164.915 138.470 167.075 ;
        RECT 140.130 164.915 153.250 167.075 ;
        RECT 81.010 150.495 86.740 156.475 ;
        RECT 88.400 150.495 94.130 156.475 ;
        RECT 95.790 150.495 101.520 156.475 ;
        RECT 103.180 150.495 108.910 156.475 ;
        RECT 110.570 150.495 116.300 156.475 ;
        RECT 117.960 150.495 123.690 156.475 ;
        RECT 125.350 150.495 131.080 156.475 ;
        RECT 132.740 150.495 138.470 156.475 ;
        RECT 140.130 150.495 145.860 156.475 ;
        RECT 147.520 150.495 153.250 156.475 ;
        RECT 81.010 136.075 86.740 142.055 ;
        RECT 88.400 136.075 94.130 142.055 ;
        RECT 95.790 136.075 101.520 142.055 ;
        RECT 103.180 136.075 108.910 142.055 ;
        RECT 110.570 136.075 116.300 142.055 ;
        RECT 117.960 136.075 123.690 142.055 ;
        RECT 125.350 136.075 131.080 142.055 ;
        RECT 132.740 136.075 138.470 142.055 ;
        RECT 140.130 136.075 145.860 142.055 ;
        RECT 147.520 136.075 153.250 142.055 ;
        RECT 81.010 121.655 86.740 127.635 ;
        RECT 88.400 121.655 94.130 127.635 ;
        RECT 95.790 121.655 101.520 127.635 ;
        RECT 103.180 121.655 108.910 127.635 ;
        RECT 110.570 121.655 116.300 127.635 ;
        RECT 117.960 121.655 123.690 127.635 ;
        RECT 125.350 121.655 131.080 127.635 ;
        RECT 132.740 121.655 138.470 127.635 ;
        RECT 140.130 121.655 145.860 127.635 ;
        RECT 147.520 121.655 153.250 127.635 ;
        RECT 6.960 107.600 20.080 109.760 ;
        RECT 21.740 107.600 34.860 109.760 ;
        RECT 36.520 107.600 49.640 109.760 ;
        RECT 51.300 107.600 64.420 109.760 ;
        RECT 66.080 107.600 79.200 109.760 ;
        RECT 81.010 107.235 86.740 113.215 ;
        RECT 88.400 107.235 94.130 113.215 ;
        RECT 95.790 107.235 101.520 113.215 ;
        RECT 103.180 107.235 108.910 113.215 ;
        RECT 110.570 107.235 116.300 113.215 ;
        RECT 117.960 107.235 123.690 113.215 ;
        RECT 125.350 107.235 131.080 113.215 ;
        RECT 132.740 107.235 138.470 113.215 ;
        RECT 140.130 107.235 145.860 113.215 ;
        RECT 147.520 107.235 153.250 113.215 ;
        RECT 6.960 98.910 12.690 104.890 ;
        RECT 14.350 98.910 20.080 104.890 ;
        RECT 21.740 98.910 27.470 104.890 ;
        RECT 29.130 98.910 34.860 104.890 ;
        RECT 36.520 98.910 42.250 104.890 ;
        RECT 43.910 98.910 49.640 104.890 ;
        RECT 51.300 98.910 57.030 104.890 ;
        RECT 58.690 98.910 64.420 104.890 ;
        RECT 66.080 98.910 71.810 104.890 ;
        RECT 73.470 98.910 79.200 104.890 ;
        RECT 6.960 90.220 12.690 96.200 ;
        RECT 14.350 90.220 20.080 96.200 ;
        RECT 21.740 90.220 27.470 96.200 ;
        RECT 29.130 90.220 34.860 96.200 ;
        RECT 36.520 90.220 42.250 96.200 ;
        RECT 43.910 90.220 49.640 96.200 ;
        RECT 51.300 90.220 57.030 96.200 ;
        RECT 58.690 90.220 64.420 96.200 ;
        RECT 66.080 90.220 71.810 96.200 ;
        RECT 73.470 90.220 79.200 96.200 ;
        RECT 81.010 92.815 86.740 98.795 ;
        RECT 88.400 92.815 94.130 98.795 ;
        RECT 95.790 92.815 101.520 98.795 ;
        RECT 103.180 92.815 108.910 98.795 ;
        RECT 110.570 92.815 116.300 98.795 ;
        RECT 117.960 92.815 123.690 98.795 ;
        RECT 125.350 92.815 131.080 98.795 ;
        RECT 132.740 92.815 138.470 98.795 ;
        RECT 140.130 92.815 145.860 98.795 ;
        RECT 147.520 92.815 153.250 98.795 ;
        RECT 6.960 81.530 12.690 87.510 ;
        RECT 14.350 81.530 20.080 87.510 ;
        RECT 21.740 81.530 27.470 87.510 ;
        RECT 29.130 81.530 34.860 87.510 ;
        RECT 36.520 81.530 42.250 87.510 ;
        RECT 43.910 81.530 49.640 87.510 ;
        RECT 51.300 81.530 57.030 87.510 ;
        RECT 58.690 81.530 64.420 87.510 ;
        RECT 66.080 81.530 71.810 87.510 ;
        RECT 73.470 81.530 79.200 87.510 ;
        RECT 6.960 72.840 12.690 78.820 ;
        RECT 14.350 72.840 20.080 78.820 ;
        RECT 21.740 72.840 27.470 78.820 ;
        RECT 29.130 72.840 34.860 78.820 ;
        RECT 36.520 72.840 42.250 78.820 ;
        RECT 43.910 72.840 49.640 78.820 ;
        RECT 51.300 72.840 57.030 78.820 ;
        RECT 58.690 72.840 64.420 78.820 ;
        RECT 66.080 72.840 71.810 78.820 ;
        RECT 73.470 72.840 79.200 78.820 ;
        RECT 81.010 78.395 86.740 84.375 ;
        RECT 88.400 78.395 94.130 84.375 ;
        RECT 95.790 78.395 101.520 84.375 ;
        RECT 103.180 78.395 108.910 84.375 ;
        RECT 110.570 78.395 116.300 84.375 ;
        RECT 117.960 78.395 123.690 84.375 ;
        RECT 125.350 78.395 131.080 84.375 ;
        RECT 132.740 78.395 138.470 84.375 ;
        RECT 140.130 78.395 145.860 84.375 ;
        RECT 147.520 78.395 153.250 84.375 ;
        RECT 6.960 64.150 12.690 70.130 ;
        RECT 14.350 64.150 20.080 70.130 ;
        RECT 21.740 64.150 27.470 70.130 ;
        RECT 29.130 64.150 34.860 70.130 ;
        RECT 36.520 64.150 42.250 70.130 ;
        RECT 43.910 64.150 49.640 70.130 ;
        RECT 51.300 64.150 57.030 70.130 ;
        RECT 58.690 64.150 64.420 70.130 ;
        RECT 66.080 64.150 71.810 70.130 ;
        RECT 73.470 64.150 79.200 70.130 ;
        RECT 81.010 63.975 86.740 69.955 ;
        RECT 88.400 63.975 94.130 69.955 ;
        RECT 95.790 63.975 101.520 69.955 ;
        RECT 103.180 63.975 108.910 69.955 ;
        RECT 110.570 63.975 116.300 69.955 ;
        RECT 117.960 63.975 123.690 69.955 ;
        RECT 125.350 63.975 131.080 69.955 ;
        RECT 132.740 63.975 138.470 69.955 ;
        RECT 140.130 63.975 145.860 69.955 ;
        RECT 147.520 63.975 153.250 69.955 ;
        RECT 6.960 55.460 12.690 61.440 ;
        RECT 14.350 55.460 20.080 61.440 ;
        RECT 21.740 55.460 27.470 61.440 ;
        RECT 29.130 55.460 34.860 61.440 ;
        RECT 36.520 55.460 42.250 61.440 ;
        RECT 43.910 55.460 49.640 61.440 ;
        RECT 51.300 55.460 57.030 61.440 ;
        RECT 58.690 55.460 64.420 61.440 ;
        RECT 66.080 55.460 71.810 61.440 ;
        RECT 73.470 55.460 79.200 61.440 ;
        RECT 6.960 46.770 12.690 52.750 ;
        RECT 14.350 46.770 20.080 52.750 ;
        RECT 21.740 46.770 27.470 52.750 ;
        RECT 29.130 46.770 34.860 52.750 ;
        RECT 36.520 46.770 42.250 52.750 ;
        RECT 43.910 46.770 49.640 52.750 ;
        RECT 51.300 46.770 57.030 52.750 ;
        RECT 58.690 46.770 64.420 52.750 ;
        RECT 66.080 46.770 71.810 52.750 ;
        RECT 73.470 46.770 79.200 52.750 ;
        RECT 81.010 49.555 86.740 55.535 ;
        RECT 88.400 49.555 94.130 55.535 ;
        RECT 95.790 49.555 101.520 55.535 ;
        RECT 103.180 49.555 108.910 55.535 ;
        RECT 110.570 49.555 116.300 55.535 ;
        RECT 117.960 49.555 123.690 55.535 ;
        RECT 125.350 49.555 131.080 55.535 ;
        RECT 132.740 49.555 138.470 55.535 ;
        RECT 140.130 49.555 145.860 55.535 ;
        RECT 147.520 49.555 153.250 55.535 ;
        RECT 6.960 38.080 12.690 44.060 ;
        RECT 14.350 38.080 20.080 44.060 ;
        RECT 21.740 38.080 27.470 44.060 ;
        RECT 29.130 38.080 34.860 44.060 ;
        RECT 36.520 38.080 42.250 44.060 ;
        RECT 43.910 38.080 49.640 44.060 ;
        RECT 51.300 38.080 57.030 44.060 ;
        RECT 58.690 38.080 64.420 44.060 ;
        RECT 66.080 38.080 71.810 44.060 ;
        RECT 73.470 38.080 79.200 44.060 ;
        RECT 6.960 29.390 12.690 35.370 ;
        RECT 14.350 29.390 20.080 35.370 ;
        RECT 21.740 29.390 27.470 35.370 ;
        RECT 29.130 29.390 34.860 35.370 ;
        RECT 36.520 29.390 42.250 35.370 ;
        RECT 43.910 29.390 49.640 35.370 ;
        RECT 51.300 29.390 57.030 35.370 ;
        RECT 58.690 29.390 64.420 35.370 ;
        RECT 66.080 29.390 71.810 35.370 ;
        RECT 73.470 29.390 79.200 35.370 ;
        RECT 81.010 35.135 86.740 41.115 ;
        RECT 88.400 35.135 94.130 41.115 ;
        RECT 95.790 35.135 101.520 41.115 ;
        RECT 103.180 35.135 108.910 41.115 ;
        RECT 110.570 35.135 116.300 41.115 ;
        RECT 117.960 35.135 123.690 41.115 ;
        RECT 125.350 35.135 131.080 41.115 ;
        RECT 132.740 35.135 138.470 41.115 ;
        RECT 140.130 35.135 145.860 41.115 ;
        RECT 147.520 35.135 153.250 41.115 ;
        RECT 6.980 24.580 12.670 26.625 ;
        RECT 14.350 24.520 27.470 26.680 ;
        RECT 29.130 24.520 42.250 26.680 ;
        RECT 43.910 24.520 57.030 26.680 ;
        RECT 58.690 24.520 71.810 26.680 ;
        RECT 73.490 24.580 79.180 26.625 ;
        RECT 81.030 24.595 86.720 26.640 ;
        RECT 88.400 24.535 101.520 26.695 ;
        RECT 103.180 24.535 116.300 26.695 ;
        RECT 117.960 24.535 131.080 26.695 ;
        RECT 132.740 24.535 145.860 26.695 ;
        RECT 147.540 24.595 153.230 26.640 ;
        RECT 144.855 20.550 145.175 20.595 ;
        RECT 8.660 20.170 9.040 20.550 ;
        RECT 144.420 20.320 150.040 20.550 ;
        RECT 144.855 20.275 145.175 20.320 ;
        RECT 105.595 19.680 105.915 19.725 ;
        RECT 102.795 19.450 114.635 19.680 ;
        RECT 11.590 16.410 24.710 18.570 ;
        RECT 26.370 16.410 39.490 18.570 ;
        RECT 41.150 16.410 54.270 18.570 ;
        RECT 55.930 16.410 69.050 18.570 ;
        RECT 70.710 16.410 83.830 18.570 ;
        RECT 103.525 18.355 103.755 19.450 ;
        RECT 105.595 19.405 105.915 19.450 ;
        RECT 144.900 19.225 145.130 20.275 ;
        RECT 144.900 19.150 145.370 19.225 ;
        RECT 144.900 18.995 145.415 19.150 ;
        RECT 145.095 18.830 145.415 18.995 ;
        RECT 104.045 18.560 104.505 18.790 ;
        RECT 107.005 18.560 107.465 18.790 ;
        RECT 109.965 18.560 110.425 18.790 ;
        RECT 112.925 18.560 113.385 18.790 ;
        RECT 103.525 18.125 103.995 18.355 ;
        RECT 91.455 15.740 97.145 17.785 ;
        RECT 103.765 17.355 103.995 18.125 ;
        RECT 104.555 17.585 104.785 18.355 ;
        RECT 106.725 17.585 106.955 18.355 ;
        RECT 104.555 17.355 105.275 17.585 ;
        RECT 104.115 17.150 104.435 17.195 ;
        RECT 104.045 16.920 104.505 17.150 ;
        RECT 104.115 16.875 104.435 16.920 ;
        RECT 104.160 16.095 104.390 16.875 ;
        RECT 104.115 15.775 104.435 16.095 ;
        RECT 104.160 14.915 104.390 15.775 ;
        RECT 105.045 14.985 105.275 17.355 ;
        RECT 106.235 17.355 106.955 17.585 ;
        RECT 107.515 17.585 107.745 18.355 ;
        RECT 109.685 17.735 109.915 18.355 ;
        RECT 109.640 17.585 109.960 17.735 ;
        RECT 107.515 17.415 109.960 17.585 ;
        RECT 110.475 17.585 110.705 18.355 ;
        RECT 112.645 17.735 112.875 18.355 ;
        RECT 112.600 17.585 112.920 17.735 ;
        RECT 107.515 17.355 109.915 17.415 ;
        RECT 110.475 17.355 111.195 17.585 ;
        RECT 103.795 14.685 104.755 14.915 ;
        RECT 105.000 14.665 105.320 14.985 ;
        RECT 105.045 14.525 105.275 14.665 ;
        RECT 103.515 13.755 103.745 14.525 ;
        RECT 103.275 13.525 103.745 13.755 ;
        RECT 104.805 14.295 105.275 14.525 ;
        RECT 106.235 14.525 106.465 17.355 ;
        RECT 107.075 17.150 107.395 17.195 ;
        RECT 107.005 16.920 107.670 17.150 ;
        RECT 107.075 16.875 107.670 16.920 ;
        RECT 106.840 15.985 107.160 16.305 ;
        RECT 106.885 14.985 107.115 15.985 ;
        RECT 107.440 15.850 107.670 16.875 ;
        RECT 107.395 15.530 107.715 15.850 ;
        RECT 106.840 14.915 107.160 14.985 ;
        RECT 106.755 14.685 107.715 14.915 ;
        RECT 106.840 14.665 107.160 14.685 ;
        RECT 108.005 14.525 108.235 17.355 ;
        RECT 109.195 14.525 109.425 17.355 ;
        RECT 109.760 16.920 110.425 17.150 ;
        RECT 109.760 16.305 109.990 16.920 ;
        RECT 110.965 16.740 111.195 17.355 ;
        RECT 112.155 17.415 112.920 17.585 ;
        RECT 113.435 17.585 113.665 18.355 ;
        RECT 114.110 17.585 114.430 17.630 ;
        RECT 112.155 17.355 112.875 17.415 ;
        RECT 113.435 17.355 114.430 17.585 ;
        RECT 110.920 16.420 111.240 16.740 ;
        RECT 109.715 15.985 110.035 16.305 ;
        RECT 110.270 15.530 110.590 15.850 ;
        RECT 110.315 14.915 110.545 15.530 ;
        RECT 109.715 14.685 110.675 14.915 ;
        RECT 110.965 14.525 111.195 16.420 ;
        RECT 106.235 14.295 106.705 14.525 ;
        RECT 104.805 13.525 105.035 14.295 ;
        RECT 106.475 13.525 106.705 14.295 ;
        RECT 107.765 14.465 109.665 14.525 ;
        RECT 107.765 14.295 109.710 14.465 ;
        RECT 107.765 13.525 107.995 14.295 ;
        RECT 109.390 14.145 109.710 14.295 ;
        RECT 110.725 14.295 111.195 14.525 ;
        RECT 112.155 14.525 112.385 17.355 ;
        RECT 114.110 17.310 114.430 17.355 ;
        RECT 113.315 17.150 113.635 17.195 ;
        RECT 112.925 16.920 113.635 17.150 ;
        RECT 113.315 16.875 113.635 16.920 ;
        RECT 112.675 14.685 113.635 14.915 ;
        RECT 114.110 14.525 114.430 14.570 ;
        RECT 112.155 14.465 112.625 14.525 ;
        RECT 112.155 14.295 112.670 14.465 ;
        RECT 109.435 13.525 109.665 14.145 ;
        RECT 110.725 13.525 110.955 14.295 ;
        RECT 112.350 14.145 112.670 14.295 ;
        RECT 113.685 14.295 114.430 14.525 ;
        RECT 130.095 14.390 135.785 16.435 ;
        RECT 143.145 15.255 143.465 15.575 ;
        RECT 112.395 13.525 112.625 14.145 ;
        RECT 113.685 13.525 113.915 14.295 ;
        RECT 114.110 14.250 114.430 14.295 ;
        RECT 143.190 13.950 143.420 15.255 ;
        RECT 145.140 15.225 145.370 18.830 ;
        RECT 145.930 15.620 146.160 19.225 ;
        RECT 146.720 19.150 146.950 19.225 ;
        RECT 146.675 18.830 146.995 19.150 ;
        RECT 145.885 15.300 146.205 15.620 ;
        RECT 145.930 15.225 146.160 15.300 ;
        RECT 146.720 15.225 146.950 18.830 ;
        RECT 147.510 15.620 147.740 19.225 ;
        RECT 148.300 19.150 148.530 19.225 ;
        RECT 148.255 18.830 148.575 19.150 ;
        RECT 147.465 15.300 147.785 15.620 ;
        RECT 147.510 15.225 147.740 15.300 ;
        RECT 148.300 15.225 148.530 18.830 ;
        RECT 149.090 15.620 149.320 19.225 ;
        RECT 149.045 15.455 149.365 15.620 ;
        RECT 149.045 15.300 149.560 15.455 ;
        RECT 149.090 15.225 149.560 15.300 ;
        RECT 147.905 15.020 148.135 15.050 ;
        RECT 145.420 14.790 145.880 15.020 ;
        RECT 146.210 14.790 146.670 15.020 ;
        RECT 147.000 14.790 147.460 15.020 ;
        RECT 147.790 14.790 148.250 15.020 ;
        RECT 148.580 14.790 149.040 15.020 ;
        RECT 145.535 13.950 145.765 14.790 ;
        RECT 143.145 13.630 143.465 13.950 ;
        RECT 145.490 13.905 145.810 13.950 ;
        RECT 146.325 13.905 146.555 14.790 ;
        RECT 147.115 13.905 147.345 14.790 ;
        RECT 147.905 13.905 148.135 14.790 ;
        RECT 148.695 13.905 148.925 14.790 ;
        RECT 149.330 13.950 149.560 15.225 ;
        RECT 145.490 13.675 148.925 13.905 ;
        RECT 145.490 13.630 145.810 13.675 ;
        RECT 103.275 12.475 103.505 13.525 ;
        RECT 107.075 13.365 107.395 13.410 ;
        RECT 110.035 13.365 110.355 13.410 ;
        RECT 112.675 13.365 112.995 13.385 ;
        RECT 103.795 13.135 104.755 13.365 ;
        RECT 106.755 13.135 107.715 13.365 ;
        RECT 109.715 13.135 110.675 13.365 ;
        RECT 112.675 13.135 113.635 13.365 ;
        RECT 107.075 13.090 107.395 13.135 ;
        RECT 110.035 13.090 110.355 13.135 ;
        RECT 112.675 13.065 112.995 13.135 ;
        RECT 145.535 12.785 145.765 13.630 ;
        RECT 146.325 12.785 146.555 13.675 ;
        RECT 147.115 12.785 147.345 13.675 ;
        RECT 147.905 12.785 148.135 13.675 ;
        RECT 148.695 12.785 148.925 13.675 ;
        RECT 149.285 13.630 149.605 13.950 ;
        RECT 145.420 12.555 145.880 12.785 ;
        RECT 146.210 12.555 146.670 12.785 ;
        RECT 147.000 12.555 147.460 12.785 ;
        RECT 147.790 12.555 148.250 12.785 ;
        RECT 148.580 12.555 149.040 12.785 ;
        RECT 102.795 11.785 114.635 12.475 ;
        RECT 149.330 12.395 149.560 13.630 ;
        RECT 103.275 10.735 103.505 11.785 ;
        RECT 107.075 11.125 107.395 11.170 ;
        RECT 110.035 11.125 110.355 11.170 ;
        RECT 113.315 11.125 113.635 11.190 ;
        RECT 103.795 10.895 104.755 11.125 ;
        RECT 106.755 10.895 107.715 11.125 ;
        RECT 109.715 10.895 110.675 11.125 ;
        RECT 112.675 10.895 113.635 11.125 ;
        RECT 107.075 10.850 107.395 10.895 ;
        RECT 110.035 10.850 110.355 10.895 ;
        RECT 113.315 10.870 113.635 10.895 ;
        RECT 103.275 10.505 103.745 10.735 ;
        RECT 103.515 9.735 103.745 10.505 ;
        RECT 104.805 9.965 105.035 10.735 ;
        RECT 106.475 9.965 106.705 10.735 ;
        RECT 104.805 9.735 105.275 9.965 ;
        RECT 103.795 9.345 104.755 9.575 ;
        RECT 104.115 9.070 104.435 9.345 ;
        RECT 104.160 8.610 104.390 9.070 ;
        RECT 104.115 8.290 104.435 8.610 ;
        RECT 11.610 5.870 17.300 7.915 ;
        RECT 18.980 5.810 32.100 7.970 ;
        RECT 33.760 5.810 46.880 7.970 ;
        RECT 48.540 5.810 61.660 7.970 ;
        RECT 63.320 5.810 76.440 7.970 ;
        RECT 78.120 5.870 83.810 7.915 ;
        RECT 104.160 7.340 104.390 8.290 ;
        RECT 105.045 7.615 105.275 9.735 ;
        RECT 106.235 9.735 106.705 9.965 ;
        RECT 107.765 9.965 107.995 10.735 ;
        RECT 109.435 10.115 109.665 10.735 ;
        RECT 109.390 9.965 109.710 10.115 ;
        RECT 107.765 9.795 109.710 9.965 ;
        RECT 110.725 9.965 110.955 10.735 ;
        RECT 112.395 10.115 112.625 10.735 ;
        RECT 112.350 9.965 112.670 10.115 ;
        RECT 107.765 9.735 109.665 9.795 ;
        RECT 110.725 9.735 111.195 9.965 ;
        RECT 106.235 8.615 106.465 9.735 ;
        RECT 106.755 9.345 107.715 9.575 ;
        RECT 106.210 8.295 106.530 8.615 ;
        RECT 91.455 5.145 97.145 7.190 ;
        RECT 104.045 7.110 104.505 7.340 ;
        RECT 105.000 7.295 105.320 7.615 ;
        RECT 105.045 6.905 105.275 7.295 ;
        RECT 103.765 6.135 103.995 6.905 ;
        RECT 103.525 5.905 103.995 6.135 ;
        RECT 104.555 6.675 105.275 6.905 ;
        RECT 106.235 6.905 106.465 8.295 ;
        RECT 106.885 8.275 107.115 9.345 ;
        RECT 107.395 8.410 107.715 8.730 ;
        RECT 106.840 7.955 107.160 8.275 ;
        RECT 107.440 7.340 107.670 8.410 ;
        RECT 107.005 7.110 107.670 7.340 ;
        RECT 108.005 6.905 108.235 9.735 ;
        RECT 109.195 6.905 109.425 9.735 ;
        RECT 109.715 9.345 110.675 9.575 ;
        RECT 110.315 8.730 110.545 9.345 ;
        RECT 110.270 8.410 110.590 8.730 ;
        RECT 110.965 8.570 111.195 9.735 ;
        RECT 112.155 9.795 112.670 9.965 ;
        RECT 113.685 9.965 113.915 10.735 ;
        RECT 114.110 9.965 114.430 10.010 ;
        RECT 112.155 9.735 112.625 9.795 ;
        RECT 113.685 9.735 114.430 9.965 ;
        RECT 109.715 7.955 110.035 8.275 ;
        RECT 110.920 8.250 111.240 8.570 ;
        RECT 109.760 7.340 109.990 7.955 ;
        RECT 109.760 7.110 110.425 7.340 ;
        RECT 110.965 6.905 111.195 8.250 ;
        RECT 106.235 6.675 106.955 6.905 ;
        RECT 104.555 5.905 104.785 6.675 ;
        RECT 106.725 5.905 106.955 6.675 ;
        RECT 107.515 6.845 109.915 6.905 ;
        RECT 107.515 6.675 109.960 6.845 ;
        RECT 107.515 5.905 107.745 6.675 ;
        RECT 109.640 6.525 109.960 6.675 ;
        RECT 110.475 6.675 111.195 6.905 ;
        RECT 112.155 6.905 112.385 9.735 ;
        RECT 114.110 9.690 114.430 9.735 ;
        RECT 112.675 9.345 113.635 9.575 ;
        RECT 145.140 8.790 145.370 12.395 ;
        RECT 145.930 12.320 146.160 12.395 ;
        RECT 145.885 12.000 146.205 12.320 ;
        RECT 145.095 8.625 145.415 8.790 ;
        RECT 144.900 8.470 145.415 8.625 ;
        RECT 144.900 8.395 145.370 8.470 ;
        RECT 145.930 8.395 146.160 12.000 ;
        RECT 146.720 8.790 146.950 12.395 ;
        RECT 147.510 12.320 147.740 12.395 ;
        RECT 147.465 12.000 147.785 12.320 ;
        RECT 146.675 8.470 146.995 8.790 ;
        RECT 146.720 8.395 146.950 8.470 ;
        RECT 147.510 8.395 147.740 12.000 ;
        RECT 148.300 8.790 148.530 12.395 ;
        RECT 149.090 12.320 149.560 12.395 ;
        RECT 149.045 12.165 149.560 12.320 ;
        RECT 149.045 12.000 149.365 12.165 ;
        RECT 148.255 8.470 148.575 8.790 ;
        RECT 148.300 8.395 148.530 8.470 ;
        RECT 149.090 8.395 149.320 12.000 ;
        RECT 112.675 7.340 112.995 7.385 ;
        RECT 144.900 7.345 145.130 8.395 ;
        RECT 112.675 7.110 113.385 7.340 ;
        RECT 144.420 7.115 150.040 7.345 ;
        RECT 112.675 7.065 112.995 7.110 ;
        RECT 114.110 6.905 114.430 6.950 ;
        RECT 112.155 6.845 112.875 6.905 ;
        RECT 112.155 6.675 112.920 6.845 ;
        RECT 109.685 5.905 109.915 6.525 ;
        RECT 110.475 5.905 110.705 6.675 ;
        RECT 112.600 6.525 112.920 6.675 ;
        RECT 113.435 6.675 114.430 6.905 ;
        RECT 112.645 5.905 112.875 6.525 ;
        RECT 113.435 5.905 113.665 6.675 ;
        RECT 114.110 6.630 114.430 6.675 ;
        RECT 103.525 4.810 103.755 5.905 ;
        RECT 104.045 5.470 104.505 5.700 ;
        RECT 107.005 5.470 107.465 5.700 ;
        RECT 109.965 5.470 110.425 5.700 ;
        RECT 112.925 5.470 113.385 5.700 ;
        RECT 105.595 4.810 105.915 4.855 ;
        RECT 102.795 4.580 114.635 4.810 ;
        RECT 105.595 4.535 105.915 4.580 ;
        RECT 130.095 3.795 135.785 5.840 ;
      LAYER met2 ;
        RECT 103.570 221.065 103.940 221.135 ;
        RECT 135.515 221.065 135.885 221.135 ;
        RECT 103.570 220.835 135.885 221.065 ;
        RECT 103.570 220.765 103.940 220.835 ;
        RECT 135.515 220.765 135.885 220.835 ;
        RECT 104.545 219.695 104.915 219.765 ;
        RECT 138.275 219.695 138.645 219.765 ;
        RECT 104.545 219.465 138.645 219.695 ;
        RECT 104.545 219.395 104.915 219.465 ;
        RECT 138.275 219.395 138.645 219.465 ;
        RECT 9.640 25.495 10.010 25.865 ;
        RECT 76.150 25.405 76.520 25.775 ;
        RECT 85.115 25.490 85.485 25.860 ;
        RECT 152.075 25.320 152.445 25.690 ;
        RECT 8.355 22.535 8.725 22.605 ;
        RECT 105.570 22.535 105.940 22.605 ;
        RECT 144.830 22.535 145.200 22.605 ;
        RECT 8.355 22.305 145.200 22.535 ;
        RECT 8.355 22.235 8.725 22.305 ;
        RECT 105.570 22.235 105.940 22.305 ;
        RECT 144.830 22.235 145.200 22.305 ;
        RECT 76.150 21.130 76.520 21.200 ;
        RECT 110.895 21.130 111.265 21.200 ;
        RECT 76.150 20.900 111.265 21.130 ;
        RECT 76.150 20.830 76.520 20.900 ;
        RECT 110.895 20.830 111.265 20.900 ;
        RECT 8.665 20.175 9.035 20.545 ;
        RECT 85.115 20.365 85.485 20.435 ;
        RECT 114.085 20.365 114.455 20.435 ;
        RECT 85.115 20.135 114.455 20.365 ;
        RECT 144.830 20.250 145.200 20.620 ;
        RECT 85.115 20.065 85.485 20.135 ;
        RECT 114.085 20.065 114.455 20.135 ;
        RECT 105.570 19.380 105.940 19.750 ;
        RECT 145.095 19.105 145.415 19.150 ;
        RECT 146.675 19.105 146.995 19.150 ;
        RECT 148.255 19.105 148.575 19.150 ;
        RECT 145.095 18.875 148.575 19.105 ;
        RECT 145.095 18.830 145.415 18.875 ;
        RECT 146.675 18.830 146.995 18.875 ;
        RECT 148.255 18.830 148.575 18.875 ;
        RECT 109.640 17.690 109.960 17.735 ;
        RECT 112.600 17.690 112.920 17.735 ;
        RECT 109.640 17.460 112.920 17.690 ;
        RECT 109.640 17.415 109.960 17.460 ;
        RECT 112.600 17.415 112.920 17.460 ;
        RECT 114.085 17.285 114.455 17.655 ;
        RECT 104.115 17.150 104.435 17.195 ;
        RECT 107.075 17.150 107.395 17.195 ;
        RECT 104.045 16.920 107.465 17.150 ;
        RECT 104.115 16.875 104.435 16.920 ;
        RECT 107.075 16.875 107.395 16.920 ;
        RECT 113.290 16.850 113.660 17.220 ;
        RECT 96.110 16.695 96.430 16.740 ;
        RECT 110.920 16.695 111.240 16.740 ;
        RECT 96.110 16.465 111.240 16.695 ;
        RECT 96.110 16.420 96.430 16.465 ;
        RECT 110.920 16.420 111.240 16.465 ;
        RECT 106.840 16.260 107.160 16.305 ;
        RECT 109.715 16.260 110.035 16.305 ;
        RECT 103.570 16.050 103.940 16.120 ;
        RECT 104.115 16.050 104.435 16.095 ;
        RECT 103.570 15.820 104.435 16.050 ;
        RECT 106.840 16.030 110.035 16.260 ;
        RECT 106.840 15.985 107.160 16.030 ;
        RECT 109.715 15.985 110.035 16.030 ;
        RECT 103.570 15.750 103.940 15.820 ;
        RECT 104.115 15.775 104.435 15.820 ;
        RECT 107.395 15.805 107.715 15.850 ;
        RECT 110.270 15.805 110.590 15.850 ;
        RECT 107.395 15.575 110.590 15.805 ;
        RECT 107.395 15.530 107.715 15.575 ;
        RECT 110.270 15.530 110.590 15.575 ;
        RECT 114.085 15.530 114.455 15.600 ;
        RECT 145.885 15.575 146.205 15.620 ;
        RECT 147.465 15.575 147.785 15.620 ;
        RECT 149.045 15.575 149.365 15.620 ;
        RECT 132.780 15.530 133.100 15.575 ;
        RECT 143.145 15.530 143.465 15.575 ;
        RECT 114.085 15.300 143.465 15.530 ;
        RECT 145.885 15.345 149.365 15.575 ;
        RECT 145.885 15.300 146.205 15.345 ;
        RECT 147.465 15.300 147.785 15.345 ;
        RECT 149.045 15.300 149.365 15.345 ;
        RECT 114.085 15.230 114.455 15.300 ;
        RECT 132.780 15.255 133.100 15.300 ;
        RECT 143.145 15.255 143.465 15.300 ;
        RECT 105.000 14.940 105.320 14.985 ;
        RECT 106.840 14.940 107.160 14.985 ;
        RECT 105.000 14.710 107.160 14.940 ;
        RECT 105.000 14.665 105.320 14.710 ;
        RECT 106.840 14.665 107.160 14.710 ;
        RECT 109.390 14.420 109.710 14.465 ;
        RECT 112.350 14.420 112.670 14.465 ;
        RECT 109.390 14.190 112.670 14.420 ;
        RECT 114.085 14.225 114.455 14.595 ;
        RECT 109.390 14.145 109.710 14.190 ;
        RECT 112.350 14.145 112.670 14.190 ;
        RECT 143.145 13.905 143.465 13.950 ;
        RECT 145.490 13.905 145.810 13.950 ;
        RECT 143.145 13.675 145.810 13.905 ;
        RECT 143.145 13.630 143.465 13.675 ;
        RECT 145.490 13.630 145.810 13.675 ;
        RECT 149.285 13.905 149.605 13.950 ;
        RECT 152.075 13.905 152.445 13.975 ;
        RECT 149.285 13.675 152.445 13.905 ;
        RECT 149.285 13.630 149.605 13.675 ;
        RECT 152.075 13.605 152.445 13.675 ;
        RECT 107.075 13.090 107.395 13.410 ;
        RECT 110.035 13.090 110.355 13.410 ;
        RECT 107.120 11.170 107.350 13.090 ;
        RECT 110.080 11.170 110.310 13.090 ;
        RECT 112.650 13.040 113.020 13.410 ;
        RECT 145.885 12.275 146.205 12.320 ;
        RECT 147.465 12.275 147.785 12.320 ;
        RECT 149.045 12.275 149.365 12.320 ;
        RECT 145.885 12.045 149.365 12.275 ;
        RECT 145.885 12.000 146.205 12.045 ;
        RECT 147.465 12.000 147.785 12.045 ;
        RECT 149.045 12.000 149.365 12.045 ;
        RECT 107.075 10.850 107.395 11.170 ;
        RECT 110.035 10.850 110.355 11.170 ;
        RECT 113.290 10.845 113.660 11.215 ;
        RECT 109.390 10.070 109.710 10.115 ;
        RECT 112.350 10.070 112.670 10.115 ;
        RECT 109.390 9.840 112.670 10.070 ;
        RECT 109.390 9.795 109.710 9.840 ;
        RECT 112.350 9.795 112.670 9.840 ;
        RECT 114.085 9.665 114.455 10.035 ;
        RECT 104.115 9.345 104.435 9.390 ;
        RECT 113.290 9.345 113.660 9.415 ;
        RECT 104.115 9.115 113.660 9.345 ;
        RECT 104.115 9.070 104.435 9.115 ;
        RECT 113.290 9.045 113.660 9.115 ;
        RECT 145.095 8.745 145.415 8.790 ;
        RECT 146.675 8.745 146.995 8.790 ;
        RECT 148.255 8.745 148.575 8.790 ;
        RECT 107.395 8.685 107.715 8.730 ;
        RECT 110.270 8.685 110.590 8.730 ;
        RECT 104.545 8.610 104.915 8.635 ;
        RECT 104.115 8.290 104.915 8.610 ;
        RECT 104.545 8.265 104.915 8.290 ;
        RECT 106.185 8.270 106.555 8.640 ;
        RECT 107.395 8.455 110.590 8.685 ;
        RECT 107.395 8.410 107.715 8.455 ;
        RECT 110.270 8.410 110.590 8.455 ;
        RECT 106.840 8.230 107.160 8.275 ;
        RECT 109.715 8.230 110.035 8.275 ;
        RECT 106.840 8.000 110.035 8.230 ;
        RECT 110.895 8.225 111.265 8.595 ;
        RECT 145.095 8.515 148.575 8.745 ;
        RECT 145.095 8.470 145.415 8.515 ;
        RECT 146.675 8.470 146.995 8.515 ;
        RECT 148.255 8.470 148.575 8.515 ;
        RECT 106.840 7.955 107.160 8.000 ;
        RECT 109.715 7.955 110.035 8.000 ;
        RECT 105.000 7.570 105.320 7.615 ;
        RECT 112.650 7.570 113.020 7.640 ;
        RECT 105.000 7.340 113.020 7.570 ;
        RECT 105.000 7.295 105.320 7.340 ;
        RECT 14.270 6.700 14.640 7.070 ;
        RECT 80.780 6.695 81.150 7.065 ;
        RECT 112.650 7.040 113.020 7.340 ;
        RECT 109.640 6.800 109.960 6.845 ;
        RECT 112.600 6.800 112.920 6.845 ;
        RECT 109.640 6.570 112.920 6.800 ;
        RECT 114.085 6.605 114.455 6.975 ;
        RECT 109.640 6.525 109.960 6.570 ;
        RECT 112.600 6.525 112.920 6.570 ;
        RECT 94.115 5.990 94.485 6.360 ;
        RECT 105.570 4.510 105.940 4.880 ;
        RECT 80.780 3.660 81.150 3.730 ;
        RECT 106.185 3.660 106.555 3.730 ;
        RECT 80.780 3.430 106.555 3.660 ;
        RECT 80.780 3.360 81.150 3.430 ;
        RECT 106.185 3.360 106.555 3.430 ;
        RECT 9.640 1.930 10.010 2.000 ;
        RECT 14.270 1.930 14.640 2.000 ;
        RECT 94.115 1.930 94.485 2.000 ;
        RECT 152.075 1.930 152.445 2.000 ;
        RECT 9.640 1.700 152.445 1.930 ;
        RECT 9.640 1.630 10.010 1.700 ;
        RECT 14.270 1.630 14.640 1.700 ;
        RECT 94.115 1.630 94.485 1.700 ;
        RECT 152.075 1.630 152.445 1.700 ;
      LAYER met3 ;
        RECT 135.510 224.675 135.890 225.055 ;
        RECT 135.550 221.115 135.850 224.675 ;
        RECT 138.270 224.635 138.650 225.015 ;
        RECT 103.590 220.785 103.920 221.115 ;
        RECT 135.535 220.785 135.865 221.115 ;
        RECT 9.660 25.515 9.990 25.845 ;
        RECT 1.860 22.570 2.420 22.700 ;
        RECT 8.375 22.570 8.705 22.585 ;
        RECT 1.860 22.270 8.705 22.570 ;
        RECT 1.860 22.140 2.420 22.270 ;
        RECT 8.375 22.255 8.705 22.270 ;
        RECT 4.635 20.510 5.195 20.640 ;
        RECT 8.685 20.510 9.015 20.525 ;
        RECT 4.635 20.210 9.015 20.510 ;
        RECT 4.635 20.080 5.195 20.210 ;
        RECT 8.685 20.195 9.015 20.210 ;
        RECT 9.675 1.980 9.975 25.515 ;
        RECT 76.170 25.425 76.500 25.755 ;
        RECT 85.135 25.510 85.465 25.840 ;
        RECT 76.185 21.180 76.485 25.425 ;
        RECT 76.170 20.850 76.500 21.180 ;
        RECT 85.150 20.415 85.450 25.510 ;
        RECT 85.135 20.085 85.465 20.415 ;
        RECT 103.605 16.100 103.905 220.785 ;
        RECT 138.310 219.745 138.610 224.635 ;
        RECT 104.565 219.415 104.895 219.745 ;
        RECT 138.295 219.415 138.625 219.745 ;
        RECT 103.590 15.770 103.920 16.100 ;
        RECT 104.580 8.615 104.880 219.415 ;
        RECT 152.095 25.340 152.425 25.670 ;
        RECT 105.590 22.255 105.920 22.585 ;
        RECT 144.850 22.255 145.180 22.585 ;
        RECT 105.605 19.730 105.905 22.255 ;
        RECT 110.915 20.850 111.245 21.180 ;
        RECT 105.590 19.400 105.920 19.730 ;
        RECT 104.565 8.285 104.895 8.615 ;
        RECT 14.290 6.720 14.620 7.050 ;
        RECT 14.305 1.980 14.605 6.720 ;
        RECT 80.800 6.715 81.130 7.045 ;
        RECT 80.815 3.710 81.115 6.715 ;
        RECT 94.135 6.010 94.465 6.340 ;
        RECT 80.800 3.380 81.130 3.710 ;
        RECT 94.150 1.980 94.450 6.010 ;
        RECT 105.605 4.860 105.905 19.400 ;
        RECT 106.205 8.290 106.535 8.620 ;
        RECT 110.930 8.575 111.230 20.850 ;
        RECT 144.865 20.600 145.165 22.255 ;
        RECT 114.105 20.085 114.435 20.415 ;
        RECT 144.850 20.270 145.180 20.600 ;
        RECT 114.120 17.635 114.420 20.085 ;
        RECT 114.105 17.305 114.435 17.635 ;
        RECT 113.310 16.870 113.640 17.200 ;
        RECT 112.670 13.060 113.000 13.390 ;
        RECT 105.590 4.530 105.920 4.860 ;
        RECT 106.220 3.710 106.520 8.290 ;
        RECT 110.915 8.245 111.245 8.575 ;
        RECT 112.685 7.620 112.985 13.060 ;
        RECT 113.325 11.195 113.625 16.870 ;
        RECT 114.120 15.580 114.420 17.305 ;
        RECT 114.105 15.250 114.435 15.580 ;
        RECT 114.120 14.575 114.420 15.250 ;
        RECT 114.105 14.245 114.435 14.575 ;
        RECT 113.310 10.865 113.640 11.195 ;
        RECT 113.325 9.395 113.625 10.865 ;
        RECT 114.120 10.015 114.420 14.245 ;
        RECT 152.110 13.955 152.410 25.340 ;
        RECT 152.095 13.625 152.425 13.955 ;
        RECT 114.105 9.685 114.435 10.015 ;
        RECT 113.310 9.065 113.640 9.395 ;
        RECT 112.670 7.060 113.000 7.620 ;
        RECT 114.120 6.955 114.420 9.685 ;
        RECT 114.105 6.625 114.435 6.955 ;
        RECT 106.205 3.380 106.535 3.710 ;
        RECT 9.660 1.650 9.990 1.980 ;
        RECT 14.290 1.650 14.620 1.980 ;
        RECT 94.135 1.650 94.465 1.980 ;
        RECT 132.790 1.000 133.090 5.090 ;
        RECT 152.110 1.980 152.410 13.625 ;
        RECT 152.095 1.650 152.425 1.980 ;
        RECT 152.110 1.000 152.410 1.650 ;
        RECT 132.750 0.620 133.130 1.000 ;
        RECT 152.070 0.620 152.450 1.000 ;
      LAYER met4 ;
        RECT 135.535 224.760 135.550 225.030 ;
        RECT 135.850 224.760 135.865 225.030 ;
        RECT 135.535 224.700 135.865 224.760 ;
        RECT 138.295 224.760 138.310 224.990 ;
        RECT 138.610 224.760 138.625 224.990 ;
        RECT 138.295 224.660 138.625 224.760 ;
  END
END tt_um_alexandercoabad_mixedsignal
END LIBRARY

