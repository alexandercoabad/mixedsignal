** sch_path: /foss/designs/mixedsignal/xschem/mixedsignal.sch
.subckt mixedsignal VDD GND S1 S2 VIN VOUT
*.PININFO VOUT:O VIN:I S1:I S2:I VDD:I GND:I
R1 VOUT mux_in 300k m=1
XM3 VOUT mux_in VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=20 nf=1 m=1
XM4 VOUT mux_in GND GND sky130_fd_pr__nfet_01v8 L=0.5 W=20 nf=1 m=1
R7 VOUT net3 300 m=1
x1 S1 S2 VDD GND net4 net1 mux_in net2 net3 4-to-1_analog_MUX
R8 VOUT net2 30k m=1
R9 mux_in VIN 3k m=1
* noconn VOUT
* noconn #net4
R2 VOUT net1 3k m=1
.ends

* expanding   symbol:  4-to-1_analog_MUX.sym # of pins=9
** sym_path: /foss/designs/mixedsignal/xschem/4-to-1_analog_MUX.sym
** sch_path: /foss/designs/mixedsignal/xschem/4-to-1_analog_MUX.sch
.subckt 4-to-1_analog_MUX S1 S2 VDD GND I1 I2 OUT I3 I4
*.PININFO I1:I I2:I I3:I I4:I OUT:O S1:I S2:I VDD:I GND:I
XM1 net1 S1 I1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 I1 S1bar net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 net1 S1bar I3 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 I3 S1 net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 net2 S1 I2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 I2 S1bar net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM7 net2 S1bar I4 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM8 I4 S1 net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
x1 S1 S1bar GND VDD Inverter
x2 S2 S2bar GND VDD Inverter
XM9 OUT S2 net1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM10 net1 S2bar OUT GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM11 OUT S2bar net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM12 net2 S2 OUT GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  Inverter.sym # of pins=4
** sym_path: /foss/designs/mixedsignal/xschem/Inverter.sym
** sch_path: /foss/designs/mixedsignal/xschem/Inverter.sch
.subckt Inverter Vin Vout GND VDD
*.PININFO Vout:O Vin:I VDD:I GND:I
XM1 Vout Vin VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 Vout Vin GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
.ends

.end
